package nn_parameters;
localparam DATA_WIDTH = 16;
localparam IN_SIZE_1 = 128;
localparam OUT_SIZE_1 = 64;




endpackage