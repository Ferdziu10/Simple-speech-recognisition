import nn_parameters::*;

module dense_layer_1 (
    input clk,
    input rst,
    input logic [15:0] input_vector [IN_SIZE_1-1:0],
    output logic signed [23:0] output_vector [OUT_SIZE_1-1:0]
);


    logic signed [7:0] weight_matrix [IN_SIZE_1-1:0][OUT_SIZE_1-1:0];
    logic signed [7:0] bias_vector [OUT_SIZE_1-1:0];
    logic signed [23:0] output_vector_nxt [OUT_SIZE_1-1:0];
    logic [7:0] i;
    logic [7:0] i_nxt;
    
    integer j, k;
    assign weight_matrix = {{8'hfd, 8'h04, 8'hfb, 8'hfa, 8'hf8, 8'hfc, 8'hfc, 8'h16, 8'hfe, 8'h0a, 8'h0a, 8'hfb, 8'h01, 8'hfa, 8'h08, 8'h01, 8'h0c, 8'h14, 8'hf9, 8'h00, 8'h18, 8'h05, 8'hf3, 8'h07, 8'h16, 8'hff, 8'h14, 8'h0e, 8'hf7, 8'h07, 8'h01, 8'h13, 8'hf8, 8'h0f, 8'hfd, 8'h02, 8'hf9, 8'hfc, 8'h17, 8'h0f, 8'h12, 8'hfa, 8'hfb, 8'hf7, 8'h0f, 8'hfd, 8'h0d, 8'h0f, 8'hfe, 8'h12, 8'hfd, 8'h06, 8'hff, 8'hfd, 8'hf9, 8'hfb, 8'hfd, 8'h0a, 8'hfe, 8'hfd, 8'h05, 8'h09, 8'h12, 8'h05, 8'hf8, 8'h06, 8'hf6, 8'hf9, 8'h05, 8'h02, 8'hfc, 8'h07, 8'h14, 8'h12, 8'h0e, 8'h0a, 8'h0d, 8'hfd, 8'hfc, 8'h15, 8'hff, 8'h17, 8'hfc, 8'h10, 8'h02, 8'h17, 8'hf6, 8'hfd, 8'hf8, 8'h02, 8'h02, 8'hf2, 8'h0b, 8'h10, 8'hf8, 8'h08, 8'h01, 8'hfb, 8'h03, 8'h01, 8'h04, 8'hf7, 8'h05, 8'h19, 8'hf4, 8'h00, 8'hf9, 8'h01, 8'hfd, 8'h16, 8'h00, 8'hf9, 8'h18, 8'hf8, 8'hfe, 8'h01, 8'hf9, 8'h09, 8'h14, 8'hf6, 8'h00, 8'hf6, 8'hf7, 8'hf9, 8'h0b, 8'h15, 8'h08, 8'h01},{8'hf3, 8'h07, 8'h02, 8'h14, 8'hed, 8'heb, 8'h06, 8'h0b, 8'h16, 8'h02, 8'h14, 8'h00, 8'hf3, 8'h0c, 8'hf8, 8'h02, 8'h13, 8'he9, 8'hf9, 8'h11, 8'hf7, 8'h01, 8'h06, 8'h00, 8'hf5, 8'hea, 8'h16, 8'h11, 8'hff, 8'hff, 8'hf4, 8'h02, 8'hdf, 8'h14, 8'h01, 8'he1, 8'hfe, 8'he4, 8'he9, 8'hef, 8'hfd, 8'hfb, 8'h00, 8'hfa, 8'heb, 8'h07, 8'hec, 8'hf4, 8'h0a, 8'h14, 8'h0b, 8'h09, 8'h0e, 8'hee, 8'hfa, 8'hef, 8'h08, 8'hec, 8'hfc, 8'he9, 8'hf3, 8'hed, 8'hf1, 8'h03, 8'hfb, 8'h0c, 8'he7, 8'hf9, 8'h02, 8'hed, 8'he1, 8'h1a, 8'h11, 8'h0d, 8'h0a, 8'hfb, 8'h0c, 8'h04, 8'hfc, 8'hfd, 8'hff, 8'h10, 8'hfe, 8'h13, 8'h0f, 8'hf2, 8'hf0, 8'hf8, 8'hee, 8'he4, 8'hf1, 8'hef, 8'hf2, 8'h0f, 8'h05, 8'h1c, 8'h0b, 8'hef, 8'hfd, 8'he9, 8'h0d, 8'h05, 8'he8, 8'he8, 8'hef, 8'h02, 8'hef, 8'h0b, 8'hf7, 8'h18, 8'hfc, 8'h07, 8'hee, 8'hf4, 8'h09, 8'h05, 8'he4, 8'hf6, 8'h12, 8'heb, 8'h08, 8'h0d, 8'hfb, 8'h02, 8'hf4, 8'hfa, 8'hee, 8'h03},{8'hff, 8'h19, 8'hf3, 8'h19, 8'h05, 8'hee, 8'h09, 8'heb, 8'he8, 8'heb, 8'h04, 8'hec, 8'h16, 8'hf6, 8'h03, 8'hf9, 8'hfc, 8'hf8, 8'h13, 8'h07, 8'h0d, 8'he7, 8'h04, 8'h08, 8'hfc, 8'h24, 8'h0d, 8'h0f, 8'hff, 8'hfe, 8'h0c, 8'h14, 8'h16, 8'hf1, 8'hf2, 8'hf4, 8'hfb, 8'hed, 8'h0f, 8'hfe, 8'hff, 8'h18, 8'h1e, 8'hef, 8'h07, 8'hee, 8'h07, 8'h12, 8'hf5, 8'h09, 8'h0e, 8'he2, 8'hf4, 8'hfe, 8'h02, 8'h08, 8'hf6, 8'h0b, 8'h1e, 8'h1b, 8'hf9, 8'hf1, 8'h0d, 8'h04, 8'he8, 8'h10, 8'h19, 8'h0e, 8'h05, 8'h08, 8'h00, 8'h29, 8'h0f, 8'h0b, 8'h0f, 8'h0b, 8'hf7, 8'he3, 8'hf3, 8'hfc, 8'hfc, 8'hf6, 8'h07, 8'hea, 8'heb, 8'hea, 8'hfe, 8'hf8, 8'hf4, 8'hf3, 8'h0e, 8'hf0, 8'hda, 8'he9, 8'hed, 8'hfc, 8'hf5, 8'h0e, 8'h18, 8'h0b, 8'hee, 8'hef, 8'h0c, 8'heb, 8'hf6, 8'hfe, 8'h09, 8'hfb, 8'h02, 8'hf4, 8'h1a, 8'hec, 8'h0c, 8'hfa, 8'hf6, 8'h06, 8'hfd, 8'hf5, 8'h0f, 8'h01, 8'h12, 8'he5, 8'h14, 8'he5, 8'hec, 8'hed, 8'h14, 8'hed},{8'he8, 8'hf8, 8'he9, 8'h00, 8'h00, 8'h0a, 8'h0c, 8'hf2, 8'hf2, 8'hf7, 8'hf4, 8'h00, 8'hf6, 8'hec, 8'hfc, 8'hfd, 8'hf3, 8'h14, 8'heb, 8'h0d, 8'h0f, 8'hed, 8'hdf, 8'he6, 8'hf7, 8'he9, 8'h01, 8'h12, 8'h02, 8'hed, 8'he3, 8'h03, 8'h0e, 8'h07, 8'he4, 8'hf5, 8'h10, 8'h09, 8'h10, 8'hf7, 8'h0a, 8'hf7, 8'h02, 8'hed, 8'h10, 8'h00, 8'h0d, 8'h0b, 8'h0c, 8'hfc, 8'heb, 8'h03, 8'h10, 8'he5, 8'h0c, 8'hfa, 8'h0d, 8'h13, 8'h07, 8'hee, 8'hfb, 8'hfc, 8'h04, 8'hf1, 8'hf5, 8'h1b, 8'hdc, 8'hf2, 8'h4f, 8'h17, 8'hf0, 8'h0d, 8'h00, 8'hfc, 8'hf5, 8'h09, 8'h11, 8'h00, 8'h20, 8'hea, 8'h0c, 8'hf0, 8'hf1, 8'h04, 8'h19, 8'hf4, 8'hf3, 8'hf9, 8'h12, 8'h0d, 8'h07, 8'h12, 8'hd9, 8'h14, 8'h0d, 8'h05, 8'h15, 8'h0a, 8'hfa, 8'h02, 8'h18, 8'hfb, 8'h10, 8'h04, 8'hed, 8'heb, 8'h15, 8'h12, 8'hfd, 8'hee, 8'h11, 8'h11, 8'hf2, 8'hf7, 8'h0c, 8'h23, 8'he3, 8'hed, 8'h0a, 8'hf4, 8'h09, 8'hfb, 8'hed, 8'h13, 8'h18, 8'h08, 8'h00, 8'h43},{8'h15, 8'hfd, 8'hf4, 8'h1b, 8'h11, 8'h1a, 8'h1b, 8'h09, 8'h1f, 8'h18, 8'hff, 8'h02, 8'h02, 8'h0c, 8'hed, 8'hdd, 8'h19, 8'h0f, 8'h0e, 8'h1a, 8'h05, 8'hff, 8'hf0, 8'hf8, 8'hf6, 8'hf7, 8'he9, 8'h0d, 8'h1d, 8'h0d, 8'hea, 8'hf3, 8'h08, 8'h0e, 8'hf8, 8'hfd, 8'hfb, 8'hff, 8'he7, 8'hed, 8'h0e, 8'hfe, 8'h14, 8'hfc, 8'h0a, 8'h0c, 8'hec, 8'h07, 8'hf4, 8'hfd, 8'he3, 8'hed, 8'hf4, 8'hf9, 8'h01, 8'hfa, 8'h14, 8'hf2, 8'h2b, 8'hf6, 8'hfe, 8'hea, 8'h00, 8'hfe, 8'hed, 8'h1b, 8'hec, 8'hd3, 8'h1c, 8'hf6, 8'hdc, 8'h12, 8'he9, 8'h05, 8'h03, 8'h0d, 8'hff, 8'hf0, 8'hff, 8'hfa, 8'h21, 8'hfe, 8'h00, 8'h16, 8'h21, 8'h0b, 8'hf0, 8'hf4, 8'hfe, 8'h17, 8'h09, 8'h09, 8'h15, 8'hf6, 8'heb, 8'h29, 8'h1e, 8'hfc, 8'h0f, 8'h08, 8'h26, 8'hfc, 8'h04, 8'h04, 8'h05, 8'h0c, 8'h00, 8'h23, 8'hf5, 8'h10, 8'he2, 8'hed, 8'he9, 8'h03, 8'h12, 8'h14, 8'hfd, 8'hfa, 8'h15, 8'he6, 8'he9, 8'hee, 8'h19, 8'h0b, 8'hf5, 8'h10, 8'h12, 8'hff},{8'h17, 8'hfc, 8'hf0, 8'hf2, 8'hef, 8'h08, 8'hf1, 8'hf5, 8'h11, 8'heb, 8'h17, 8'h05, 8'h12, 8'h14, 8'hea, 8'hef, 8'h03, 8'h03, 8'hfb, 8'he9, 8'hea, 8'h11, 8'hf7, 8'hdf, 8'h02, 8'h25, 8'h04, 8'hea, 8'h10, 8'h1c, 8'h08, 8'h17, 8'h05, 8'hec, 8'hf5, 8'he4, 8'hf5, 8'h03, 8'h15, 8'h0a, 8'hed, 8'hf7, 8'h03, 8'hff, 8'hf4, 8'h0e, 8'h07, 8'h0c, 8'hfd, 8'hf6, 8'h07, 8'hec, 8'hfe, 8'hd4, 8'hf3, 8'hea, 8'h16, 8'h04, 8'h11, 8'hf5, 8'hff, 8'h0e, 8'hfa, 8'he9, 8'h19, 8'hf6, 8'he5, 8'hcf, 8'he6, 8'hee, 8'he3, 8'h08, 8'h18, 8'h12, 8'h00, 8'h11, 8'hf0, 8'h01, 8'h01, 8'h07, 8'h1d, 8'h22, 8'hea, 8'hf8, 8'hdc, 8'h07, 8'hec, 8'hee, 8'h08, 8'h02, 8'h0a, 8'hed, 8'h17, 8'hff, 8'hf0, 8'hfe, 8'he7, 8'hf9, 8'hf8, 8'h06, 8'h09, 8'h1a, 8'hfa, 8'h00, 8'hf8, 8'he4, 8'hf7, 8'h0b, 8'h00, 8'h18, 8'h04, 8'hfe, 8'hf3, 8'h1b, 8'hf3, 8'hf3, 8'hf9, 8'hfa, 8'hed, 8'hed, 8'h04, 8'hf7, 8'h00, 8'hf0, 8'h06, 8'hf4, 8'hfe, 8'hf4},{8'hdc, 8'h03, 8'h17, 8'h0d, 8'h0a, 8'h0e, 8'hf3, 8'hfd, 8'h0d, 8'h06, 8'hf6, 8'hfe, 8'h10, 8'hee, 8'hf2, 8'hf4, 8'hed, 8'hee, 8'h17, 8'hf7, 8'hf6, 8'h01, 8'h09, 8'h08, 8'hff, 8'h07, 8'hea, 8'h13, 8'hea, 8'h1b, 8'h13, 8'h05, 8'h07, 8'hf9, 8'hee, 8'hef, 8'h1a, 8'hf8, 8'hf4, 8'hff, 8'hee, 8'hfd, 8'hf4, 8'h06, 8'h13, 8'h07, 8'hef, 8'h05, 8'h05, 8'h02, 8'hfe, 8'h1d, 8'h08, 8'h10, 8'h00, 8'hd7, 8'hee, 8'hfb, 8'hc4, 8'hf1, 8'h14, 8'hf4, 8'h09, 8'h03, 8'h03, 8'h06, 8'h01, 8'hef, 8'had, 8'hf3, 8'hf7, 8'h0f, 8'hf4, 8'hef, 8'h18, 8'hff, 8'hff, 8'h24, 8'hd8, 8'h14, 8'h1d, 8'h0a, 8'h00, 8'h0a, 8'h06, 8'hea, 8'h0f, 8'hfb, 8'h03, 8'he9, 8'h17, 8'hf9, 8'h25, 8'hfd, 8'hf2, 8'hfd, 8'h0d, 8'hf6, 8'hee, 8'h0e, 8'hd4, 8'hed, 8'h14, 8'heb, 8'hf1, 8'hf3, 8'he7, 8'hbe, 8'heb, 8'h08, 8'h0c, 8'h09, 8'h04, 8'he1, 8'h0d, 8'he4, 8'h1b, 8'h2c, 8'he9, 8'h0e, 8'hf1, 8'hed, 8'h0c, 8'h14, 8'hf8, 8'h02, 8'h09, 8'hf6},{8'h07, 8'h0a, 8'h07, 8'h0c, 8'hdf, 8'he3, 8'hef, 8'h12, 8'hf9, 8'hf0, 8'hf3, 8'h11, 8'he0, 8'he1, 8'hf7, 8'hf4, 8'h19, 8'h0b, 8'h0e, 8'hf4, 8'h05, 8'h00, 8'hf9, 8'h15, 8'h0c, 8'hdc, 8'hf3, 8'h19, 8'h06, 8'h07, 8'h36, 8'h00, 8'h10, 8'h0d, 8'h0e, 8'he2, 8'h04, 8'hf2, 8'h03, 8'h14, 8'h01, 8'hf8, 8'h2e, 8'h0d, 8'hfa, 8'hfc, 8'hf5, 8'hf0, 8'hdd, 8'h16, 8'h1d, 8'hfe, 8'h09, 8'h1a, 8'h09, 8'h1f, 8'hff, 8'h2a, 8'h2d, 8'h13, 8'hf4, 8'h10, 8'hf9, 8'h09, 8'h1b, 8'hf9, 8'hf7, 8'hf1, 8'he8, 8'h16, 8'h13, 8'h08, 8'hf5, 8'hfc, 8'hf8, 8'h20, 8'h08, 8'hfc, 8'hed, 8'h04, 8'hd0, 8'h12, 8'hee, 8'h07, 8'hc8, 8'hfa, 8'h08, 8'heb, 8'he8, 8'h0d, 8'hf8, 8'hfe, 8'h1e, 8'h12, 8'h0d, 8'hf9, 8'hf4, 8'h0c, 8'h05, 8'hfb, 8'hea, 8'hec, 8'h01, 8'hea, 8'hdd, 8'h1f, 8'hec, 8'h0c, 8'h0e, 8'hf7, 8'hea, 8'h11, 8'h06, 8'hf5, 8'h0b, 8'hee, 8'h20, 8'he9, 8'h14, 8'h11, 8'hfa, 8'hee, 8'he4, 8'hde, 8'h04, 8'h02, 8'h10, 8'hd8},{8'hf8, 8'hea, 8'h23, 8'he6, 8'hf6, 8'h0f, 8'h1a, 8'h19, 8'hfc, 8'h01, 8'h03, 8'h03, 8'hdd, 8'h12, 8'h11, 8'he7, 8'h09, 8'hfb, 8'hff, 8'he4, 8'h0b, 8'hf9, 8'hf1, 8'hf1, 8'hf1, 8'h11, 8'h09, 8'hee, 8'hed, 8'hf3, 8'heb, 8'h00, 8'hfc, 8'heb, 8'hf4, 8'hd4, 8'hff, 8'h03, 8'h06, 8'hfc, 8'h0d, 8'hf3, 8'h07, 8'h16, 8'hf9, 8'he4, 8'h03, 8'hf0, 8'h01, 8'hfa, 8'h03, 8'h1b, 8'h06, 8'h1e, 8'hee, 8'h04, 8'h20, 8'hcd, 8'h07, 8'hfe, 8'hfe, 8'hfa, 8'hfa, 8'hf9, 8'h17, 8'h1d, 8'hf7, 8'heb, 8'hde, 8'h00, 8'h13, 8'h08, 8'h0d, 8'hf1, 8'h03, 8'h17, 8'h08, 8'h3a, 8'hd7, 8'hf1, 8'h38, 8'h09, 8'h06, 8'h04, 8'h13, 8'h02, 8'h00, 8'hea, 8'hfd, 8'hce, 8'h10, 8'h0b, 8'h2c, 8'h13, 8'he8, 8'h1a, 8'hd1, 8'h0f, 8'he8, 8'h0c, 8'hfb, 8'he6, 8'h16, 8'h0e, 8'hff, 8'he2, 8'h0d, 8'h03, 8'hf6, 8'h03, 8'hcc, 8'hfd, 8'h02, 8'h12, 8'h0c, 8'hfb, 8'h03, 8'h16, 8'h05, 8'hf0, 8'hfb, 8'h06, 8'h0c, 8'h05, 8'h00, 8'h13, 8'h07, 8'hf0},{8'h21, 8'hf4, 8'hee, 8'h00, 8'he3, 8'hdd, 8'hff, 8'h10, 8'h16, 8'h01, 8'hed, 8'hf1, 8'hf6, 8'h03, 8'hf4, 8'h03, 8'hf7, 8'h14, 8'h0a, 8'hff, 8'hf0, 8'hfd, 8'hfd, 8'h01, 8'h18, 8'hea, 8'hf5, 8'h07, 8'h00, 8'h00, 8'h09, 8'he8, 8'hf4, 8'hf2, 8'hed, 8'h02, 8'hea, 8'h0f, 8'hef, 8'h12, 8'h19, 8'hf4, 8'he9, 8'h17, 8'h07, 8'h1d, 8'heb, 8'hf9, 8'h07, 8'h07, 8'h03, 8'hf3, 8'hdc, 8'h1f, 8'h18, 8'h07, 8'he6, 8'h32, 8'hf4, 8'hfb, 8'h02, 8'h0d, 8'h07, 8'h10, 8'hf4, 8'he1, 8'h0d, 8'h14, 8'he3, 8'he9, 8'h0c, 8'hfc, 8'h0b, 8'hf6, 8'hff, 8'hf9, 8'hef, 8'hd7, 8'h25, 8'h0e, 8'hd3, 8'hfc, 8'h00, 8'heb, 8'hf6, 8'hf5, 8'h0f, 8'hf8, 8'h1e, 8'hf4, 8'hf4, 8'h1c, 8'h09, 8'hfa, 8'h14, 8'he7, 8'h12, 8'h00, 8'h0b, 8'hfd, 8'hd2, 8'h13, 8'he7, 8'h18, 8'hfd, 8'h26, 8'hea, 8'h07, 8'hfa, 8'h13, 8'h17, 8'he9, 8'hf3, 8'hfb, 8'hf1, 8'he9, 8'h11, 8'h1a, 8'hfa, 8'h1b, 8'h14, 8'he3, 8'hdc, 8'he9, 8'h01, 8'h16, 8'h05, 8'h17},{8'h27, 8'h0f, 8'h00, 8'h11, 8'he6, 8'hee, 8'hef, 8'hf4, 8'h1a, 8'h0f, 8'h03, 8'h20, 8'h28, 8'hfc, 8'h11, 8'hf1, 8'hf5, 8'he9, 8'hea, 8'h1d, 8'hef, 8'h12, 8'h2d, 8'h0a, 8'hf3, 8'hfe, 8'heb, 8'h0c, 8'hf6, 8'hea, 8'h1a, 8'h02, 8'h11, 8'h05, 8'h14, 8'h15, 8'he6, 8'h08, 8'hf0, 8'hf0, 8'h0d, 8'h0b, 8'hf8, 8'hf0, 8'hee, 8'h0d, 8'hfe, 8'h00, 8'he5, 8'hec, 8'h02, 8'hed, 8'hf2, 8'h07, 8'h0e, 8'h1e, 8'hf6, 8'hec, 8'h0c, 8'h09, 8'h0d, 8'h00, 8'hef, 8'heb, 8'hf7, 8'h02, 8'h00, 8'h05, 8'h1a, 8'h0c, 8'h14, 8'hf1, 8'he8, 8'hf9, 8'h0b, 8'h18, 8'hfc, 8'hda, 8'h1c, 8'h12, 8'he2, 8'hf1, 8'h11, 8'heb, 8'h00, 8'h0f, 8'h13, 8'h04, 8'hff, 8'h06, 8'h06, 8'hf9, 8'h36, 8'h0b, 8'h05, 8'hf7, 8'hf8, 8'hfd, 8'hf4, 8'hfc, 8'h05, 8'hf0, 8'hf2, 8'h12, 8'hdd, 8'h0a, 8'h06, 8'h03, 8'h03, 8'hec, 8'h37, 8'hf4, 8'h16, 8'hff, 8'h0c, 8'hf2, 8'hf4, 8'he5, 8'hf7, 8'h22, 8'hfb, 8'h04, 8'hef, 8'heb, 8'hf2, 8'h01, 8'hef, 8'hef},{8'h0e, 8'hec, 8'h17, 8'h03, 8'h20, 8'h03, 8'h0a, 8'hee, 8'hde, 8'h0c, 8'hf9, 8'he2, 8'h14, 8'he3, 8'heb, 8'h16, 8'h0a, 8'h09, 8'hff, 8'hfc, 8'h10, 8'h04, 8'h0a, 8'hf3, 8'h0c, 8'h1c, 8'h08, 8'h08, 8'hdb, 8'hf1, 8'h37, 8'hfd, 8'hfb, 8'h10, 8'h04, 8'hff, 8'h13, 8'hf8, 8'h15, 8'h16, 8'hff, 8'hed, 8'hff, 8'h01, 8'hf8, 8'hf9, 8'hfc, 8'h17, 8'h10, 8'hfd, 8'h17, 8'h31, 8'h0b, 8'h12, 8'hfd, 8'h08, 8'hf9, 8'h16, 8'hef, 8'h2d, 8'hf3, 8'hea, 8'hf0, 8'h0b, 8'hf9, 8'hda, 8'h1a, 8'h02, 8'hee, 8'h14, 8'h26, 8'hfe, 8'h18, 8'hed, 8'hf6, 8'hf3, 8'hf8, 8'h1b, 8'hce, 8'h01, 8'h04, 8'hef, 8'h0d, 8'hf0, 8'he1, 8'he8, 8'h0c, 8'hf6, 8'hde, 8'hbc, 8'h1f, 8'hed, 8'hf8, 8'h08, 8'h03, 8'hfe, 8'heb, 8'h18, 8'hf4, 8'h08, 8'hcc, 8'hf3, 8'hff, 8'hff, 8'hf2, 8'h15, 8'hf8, 8'hf3, 8'h07, 8'hfe, 8'h04, 8'hfb, 8'hf5, 8'hf2, 8'h0e, 8'he9, 8'h0c, 8'h0c, 8'h14, 8'h10, 8'h19, 8'hf1, 8'h1e, 8'hdd, 8'hec, 8'hef, 8'hf0, 8'hfa},{8'h01, 8'h05, 8'hf1, 8'h02, 8'h11, 8'h13, 8'h02, 8'h19, 8'h26, 8'hfe, 8'hfd, 8'h0b, 8'h32, 8'hea, 8'h05, 8'h0a, 8'h07, 8'hf2, 8'h17, 8'hea, 8'h12, 8'h0e, 8'h04, 8'h0f, 8'h04, 8'h32, 8'hf5, 8'hee, 8'he4, 8'h2c, 8'h1c, 8'h0a, 8'h22, 8'he8, 8'hfe, 8'h03, 8'h08, 8'h08, 8'h17, 8'h06, 8'h0f, 8'hee, 8'hf6, 8'hf7, 8'hf0, 8'hee, 8'h13, 8'h10, 8'h20, 8'h0a, 8'h09, 8'he7, 8'hf6, 8'h02, 8'h15, 8'hf0, 8'h12, 8'hf9, 8'hd5, 8'h0f, 8'h11, 8'he5, 8'h04, 8'h10, 8'h1e, 8'hde, 8'h25, 8'h03, 8'he9, 8'h0e, 8'h2c, 8'hf4, 8'h03, 8'h08, 8'h09, 8'h00, 8'hfa, 8'h12, 8'hf0, 8'hef, 8'h0c, 8'h1f, 8'hff, 8'hf3, 8'hde, 8'h0b, 8'hff, 8'hfd, 8'hfd, 8'h10, 8'h33, 8'h17, 8'hf9, 8'hfd, 8'h28, 8'h09, 8'h23, 8'hef, 8'he8, 8'he9, 8'hd7, 8'hfe, 8'h07, 8'he8, 8'h00, 8'h18, 8'he9, 8'h07, 8'hf9, 8'h0a, 8'h22, 8'hf1, 8'hf6, 8'h0c, 8'he9, 8'hed, 8'h20, 8'h11, 8'h04, 8'h28, 8'h13, 8'hf8, 8'hf6, 8'h08, 8'h18, 8'hf2, 8'h08, 8'h26},{8'h08, 8'he8, 8'hff, 8'he9, 8'hfe, 8'hfc, 8'heb, 8'h17, 8'hf0, 8'hf2, 8'hfc, 8'hff, 8'h0e, 8'he7, 8'hfd, 8'hf4, 8'he8, 8'h07, 8'hfc, 8'h01, 8'h0a, 8'hef, 8'hea, 8'h10, 8'h01, 8'h0b, 8'hf7, 8'h0c, 8'he3, 8'h07, 8'h08, 8'h04, 8'h06, 8'hf5, 8'hfc, 8'h0d, 8'h05, 8'hfb, 8'h05, 8'hf6, 8'h0d, 8'he9, 8'hdd, 8'h0b, 8'h0c, 8'h04, 8'h07, 8'h05, 8'hf0, 8'hea, 8'hf2, 8'h09, 8'he8, 8'h05, 8'h00, 8'hff, 8'hed, 8'h0c, 8'hd5, 8'h08, 8'hf8, 8'h19, 8'h09, 8'h04, 8'h05, 8'h01, 8'h00, 8'hf3, 8'hfe, 8'hef, 8'h03, 8'hf6, 8'hf3, 8'he7, 8'hee, 8'h12, 8'hf0, 8'hfa, 8'hf3, 8'h02, 8'hfb, 8'h0c, 8'hfc, 8'hf3, 8'h14, 8'hfe, 8'h09, 8'h04, 8'hfd, 8'h13, 8'h11, 8'he1, 8'h17, 8'hed, 8'he5, 8'hea, 8'h0b, 8'hfa, 8'he8, 8'hf5, 8'h12, 8'hed, 8'he8, 8'hed, 8'hf2, 8'h0b, 8'he9, 8'hf7, 8'h0f, 8'hf6, 8'h04, 8'heb, 8'h04, 8'hf5, 8'h01, 8'hed, 8'h0b, 8'h15, 8'h13, 8'hf6, 8'h0e, 8'he5, 8'he3, 8'he6, 8'hfc, 8'hee, 8'hed, 8'hf3},{8'h05, 8'hf2, 8'hfd, 8'hf9, 8'he9, 8'h12, 8'hf8, 8'h0c, 8'hee, 8'hf8, 8'hec, 8'h0a, 8'hed, 8'hf9, 8'h0b, 8'h0b, 8'hef, 8'h06, 8'hfd, 8'hf1, 8'h04, 8'h05, 8'he1, 8'h0a, 8'h16, 8'he9, 8'hf6, 8'h02, 8'heb, 8'hef, 8'hf2, 8'h04, 8'hf5, 8'h17, 8'hed, 8'h0d, 8'heb, 8'hf8, 8'h09, 8'h04, 8'hea, 8'hf1, 8'h00, 8'hfc, 8'hf9, 8'he7, 8'hfa, 8'h0c, 8'h05, 8'hee, 8'he1, 8'heb, 8'h09, 8'h03, 8'he8, 8'hea, 8'h11, 8'h00, 8'h07, 8'hfe, 8'h00, 8'hf5, 8'heb, 8'hf9, 8'h00, 8'h1a, 8'hfa, 8'hee, 8'h05, 8'h0e, 8'h02, 8'hf0, 8'h15, 8'hef, 8'he8, 8'h0d, 8'h12, 8'h1a, 8'hf7, 8'h0e, 8'h13, 8'he3, 8'h0f, 8'h00, 8'he6, 8'h17, 8'hef, 8'hfe, 8'hf3, 8'hf0, 8'hee, 8'hf4, 8'hec, 8'h13, 8'h06, 8'h0c, 8'he7, 8'he7, 8'hea, 8'hf8, 8'h06, 8'hf3, 8'hf3, 8'hee, 8'hea, 8'hfe, 8'hfe, 8'hf6, 8'he6, 8'hf4, 8'hec, 8'h0d, 8'h13, 8'hfb, 8'hfe, 8'h00, 8'he7, 8'hfb, 8'he9, 8'h02, 8'hf6, 8'he5, 8'h01, 8'h0a, 8'h14, 8'hf9, 8'h00, 8'hf6},{8'h11, 8'h0e, 8'hf4, 8'hf6, 8'h05, 8'h03, 8'h0c, 8'hfc, 8'h12, 8'hf5, 8'hee, 8'hdc, 8'hf8, 8'h08, 8'h07, 8'h0d, 8'h0b, 8'h0a, 8'h00, 8'hf1, 8'h07, 8'hf4, 8'h03, 8'h0a, 8'h03, 8'h09, 8'hf4, 8'he7, 8'h14, 8'he8, 8'he6, 8'h13, 8'h08, 8'hee, 8'h0b, 8'h12, 8'heb, 8'h12, 8'hf4, 8'h14, 8'he8, 8'h03, 8'h18, 8'hdd, 8'h0c, 8'hf0, 8'h06, 8'he8, 8'h0a, 8'hf5, 8'hf3, 8'h09, 8'h0d, 8'hf6, 8'h02, 8'h12, 8'hd8, 8'hee, 8'h3b, 8'hfa, 8'hf0, 8'h08, 8'h17, 8'h00, 8'hdb, 8'h0c, 8'he7, 8'hf4, 8'hf3, 8'h0e, 8'he7, 8'h05, 8'hfb, 8'h13, 8'h00, 8'he4, 8'hf1, 8'hf1, 8'h1b, 8'hec, 8'he7, 8'h0c, 8'hf0, 8'h05, 8'h01, 8'h05, 8'he9, 8'hf9, 8'hf2, 8'h04, 8'hee, 8'hfe, 8'h09, 8'hec, 8'h05, 8'h13, 8'h0d, 8'he6, 8'h01, 8'h12, 8'hd8, 8'he8, 8'hf4, 8'hfa, 8'h03, 8'hfa, 8'h02, 8'h0f, 8'h07, 8'h02, 8'hf7, 8'he1, 8'h05, 8'h03, 8'hf8, 8'h0f, 8'hdb, 8'h15, 8'h11, 8'h02, 8'he9, 8'h02, 8'hec, 8'hf8, 8'hec, 8'hfc, 8'h0c, 8'h16},{8'hf7, 8'hed, 8'hf1, 8'hf7, 8'he0, 8'h07, 8'h11, 8'hf8, 8'hec, 8'hfa, 8'he8, 8'hff, 8'he1, 8'hff, 8'hf3, 8'h00, 8'h10, 8'h03, 8'hf3, 8'h02, 8'heb, 8'hfb, 8'hef, 8'h13, 8'h0a, 8'hed, 8'hfb, 8'hfa, 8'hfc, 8'hea, 8'h08, 8'he9, 8'he5, 8'hed, 8'hf1, 8'hf0, 8'h07, 8'he7, 8'hf2, 8'hee, 8'h0c, 8'h0c, 8'hf1, 8'hfd, 8'h06, 8'hf8, 8'hef, 8'h0a, 8'hfc, 8'hf3, 8'hfd, 8'h0f, 8'he9, 8'he9, 8'h0c, 8'h0e, 8'hef, 8'h17, 8'hfe, 8'h0c, 8'hf3, 8'h04, 8'h05, 8'hfb, 8'h02, 8'h01, 8'hf4, 8'h00, 8'h2f, 8'hf6, 8'he4, 8'hfb, 8'h09, 8'h17, 8'h0d, 8'hec, 8'h07, 8'he8, 8'h1f, 8'hfe, 8'he7, 8'heb, 8'he5, 8'he8, 8'hfc, 8'h10, 8'hf7, 8'h0f, 8'h15, 8'h22, 8'hed, 8'h08, 8'h0d, 8'hf8, 8'hed, 8'h05, 8'h0d, 8'h15, 8'hfe, 8'h0d, 8'h0f, 8'h00, 8'he9, 8'h01, 8'hd6, 8'hff, 8'h02, 8'heb, 8'he4, 8'he9, 8'h19, 8'hf9, 8'hf1, 8'hfe, 8'hf7, 8'h0f, 8'he6, 8'h15, 8'h03, 8'h07, 8'he5, 8'he0, 8'heb, 8'hf0, 8'hee, 8'hf6, 8'h11, 8'h12},{8'he9, 8'hfc, 8'h03, 8'hff, 8'he8, 8'h08, 8'hfa, 8'hf6, 8'hf7, 8'h11, 8'hfe, 8'h07, 8'heb, 8'hfa, 8'hfc, 8'hff, 8'h0f, 8'hee, 8'he4, 8'hfc, 8'h19, 8'he8, 8'hf9, 8'h03, 8'hf6, 8'he4, 8'hfb, 8'hef, 8'hf7, 8'h22, 8'h1f, 8'h0b, 8'hff, 8'h0e, 8'h03, 8'hfc, 8'hf5, 8'hf6, 8'h04, 8'hf0, 8'hff, 8'hf4, 8'h03, 8'hdf, 8'h12, 8'h00, 8'h15, 8'h12, 8'hff, 8'h05, 8'h06, 8'hfd, 8'h0e, 8'h04, 8'he0, 8'h04, 8'h07, 8'h09, 8'h01, 8'hef, 8'h18, 8'h11, 8'hfc, 8'hec, 8'hea, 8'h05, 8'hf4, 8'h02, 8'he8, 8'h16, 8'h0e, 8'h00, 8'h16, 8'h0f, 8'h02, 8'hfb, 8'h0e, 8'h01, 8'he7, 8'h10, 8'he8, 8'h09, 8'hea, 8'hf8, 8'hf2, 8'h03, 8'hea, 8'hdd, 8'hf3, 8'hf0, 8'h05, 8'h12, 8'h02, 8'h0f, 8'hf0, 8'hfc, 8'hdf, 8'h0f, 8'hea, 8'h06, 8'he7, 8'he5, 8'hf1, 8'h09, 8'hec, 8'he4, 8'h06, 8'hf8, 8'h0d, 8'h14, 8'hec, 8'hf3, 8'h14, 8'hf5, 8'he6, 8'h0c, 8'h02, 8'h25, 8'he7, 8'hec, 8'he8, 8'h09, 8'he5, 8'hef, 8'h19, 8'h0c, 8'hf7, 8'hf0},{8'hf9, 8'hfa, 8'he9, 8'hec, 8'hf1, 8'hef, 8'hfc, 8'hf6, 8'hfe, 8'hfe, 8'h02, 8'he9, 8'h1c, 8'hf9, 8'hf3, 8'heb, 8'h11, 8'h02, 8'he9, 8'h0d, 8'he9, 8'hf0, 8'hd9, 8'hee, 8'h0a, 8'h19, 8'hf9, 8'h0b, 8'h01, 8'h02, 8'h28, 8'h02, 8'heb, 8'hf9, 8'h1d, 8'hfb, 8'hfc, 8'h18, 8'hef, 8'h09, 8'hfa, 8'hf4, 8'hfe, 8'hfe, 8'hf5, 8'hfb, 8'hfe, 8'h0b, 8'h0b, 8'h05, 8'he6, 8'h12, 8'h0d, 8'h15, 8'hea, 8'he1, 8'h10, 8'h05, 8'he7, 8'hea, 8'h0f, 8'hf7, 8'hf2, 8'h05, 8'he8, 8'he3, 8'he4, 8'hea, 8'h06, 8'h12, 8'h12, 8'hf1, 8'h0c, 8'h13, 8'h18, 8'h18, 8'h11, 8'hf4, 8'hf5, 8'hf1, 8'h12, 8'h09, 8'h02, 8'hf8, 8'hef, 8'h00, 8'hed, 8'hf8, 8'hfb, 8'hfa, 8'h17, 8'hec, 8'hf9, 8'hf6, 8'hf7, 8'h0a, 8'h14, 8'h07, 8'hf1, 8'hfc, 8'hef, 8'h04, 8'h02, 8'h12, 8'h0c, 8'h0e, 8'h07, 8'hf9, 8'hf0, 8'h08, 8'h15, 8'hf7, 8'h14, 8'h00, 8'hdf, 8'hf3, 8'hee, 8'h0b, 8'h12, 8'hef, 8'h06, 8'hef, 8'h0f, 8'h04, 8'hfb, 8'h13, 8'hf7, 8'h0c},{8'hfe, 8'h08, 8'hde, 8'hea, 8'h10, 8'hf1, 8'hec, 8'h09, 8'h15, 8'hf6, 8'he8, 8'he7, 8'h1c, 8'he7, 8'heb, 8'hfa, 8'he9, 8'hf0, 8'hee, 8'hea, 8'h10, 8'he8, 8'hfb, 8'h05, 8'hf0, 8'h2a, 8'h0b, 8'hea, 8'hfc, 8'h1a, 8'h30, 8'hfa, 8'h0b, 8'he7, 8'h0f, 8'hf1, 8'hdd, 8'h21, 8'hf6, 8'h14, 8'hf4, 8'h0f, 8'h0e, 8'hdb, 8'hf4, 8'hf7, 8'hf3, 8'hed, 8'hed, 8'h06, 8'h09, 8'hf0, 8'h07, 8'h17, 8'h0a, 8'h10, 8'h0f, 8'h1d, 8'hfa, 8'h11, 8'h05, 8'hea, 8'hec, 8'h0c, 8'h03, 8'h0d, 8'h09, 8'h19, 8'hef, 8'h00, 8'h19, 8'hfe, 8'hff, 8'h09, 8'h12, 8'h0f, 8'h12, 8'he3, 8'hfe, 8'hed, 8'h09, 8'hf0, 8'h0c, 8'h16, 8'hec, 8'hfb, 8'hf3, 8'he5, 8'he7, 8'hea, 8'h2b, 8'hec, 8'h09, 8'h0e, 8'hfb, 8'h17, 8'hf8, 8'h02, 8'h15, 8'h11, 8'hea, 8'hfe, 8'h04, 8'hec, 8'hf1, 8'h05, 8'hf8, 8'h05, 8'hf8, 8'he8, 8'h14, 8'hf5, 8'h0a, 8'hf7, 8'h03, 8'h0c, 8'hf2, 8'he9, 8'hf2, 8'hff, 8'he7, 8'he3, 8'h0f, 8'hf4, 8'h16, 8'he8, 8'h0b, 8'h01},{8'he9, 8'hed, 8'he4, 8'hfa, 8'hfc, 8'hfb, 8'h09, 8'heb, 8'h05, 8'hec, 8'hfb, 8'hed, 8'h1b, 8'h09, 8'hff, 8'h0d, 8'h07, 8'h03, 8'h04, 8'h03, 8'h0e, 8'hfe, 8'hf1, 8'hfb, 8'h11, 8'h1b, 8'h11, 8'h08, 8'h0e, 8'h0a, 8'hf7, 8'h18, 8'he8, 8'h0f, 8'h16, 8'hf7, 8'hfc, 8'h14, 8'hf9, 8'he7, 8'hf2, 8'hea, 8'h02, 8'he3, 8'h03, 8'hf0, 8'he8, 8'h0e, 8'hee, 8'h14, 8'hfd, 8'hf9, 8'h02, 8'hff, 8'h0a, 8'he9, 8'hfa, 8'h12, 8'h06, 8'h11, 8'hef, 8'hfd, 8'h03, 8'hf5, 8'hd6, 8'hea, 8'h06, 8'hff, 8'h11, 8'hf4, 8'h0a, 8'h06, 8'h16, 8'h0b, 8'hf2, 8'hfd, 8'hee, 8'he4, 8'hf7, 8'h08, 8'hfa, 8'h06, 8'h06, 8'h12, 8'hfc, 8'h14, 8'he3, 8'h04, 8'h05, 8'hf0, 8'h10, 8'he7, 8'h08, 8'h01, 8'h0e, 8'h1c, 8'h0b, 8'h05, 8'h0c, 8'hf6, 8'heb, 8'hfe, 8'hf8, 8'hfc, 8'hdf, 8'h11, 8'hef, 8'h11, 8'hfd, 8'hf0, 8'h17, 8'hed, 8'hf6, 8'he9, 8'h05, 8'h0f, 8'h01, 8'hfd, 8'hf5, 8'h06, 8'h07, 8'hf6, 8'hdc, 8'hf7, 8'h14, 8'h01, 8'heb, 8'h1d},{8'h09, 8'h13, 8'h10, 8'hf0, 8'hfc, 8'hf2, 8'hf4, 8'hf5, 8'h10, 8'h06, 8'h00, 8'h00, 8'h2a, 8'h05, 8'h00, 8'he5, 8'hed, 8'hed, 8'h07, 8'hf7, 8'h0f, 8'hfa, 8'hf3, 8'he7, 8'hef, 8'h05, 8'h19, 8'hea, 8'hdf, 8'h0b, 8'h0e, 8'h0f, 8'he5, 8'hfa, 8'hf3, 8'hfa, 8'hef, 8'h12, 8'h02, 8'h05, 8'hea, 8'h0f, 8'hef, 8'hf2, 8'h0b, 8'h07, 8'h07, 8'h01, 8'h11, 8'hf0, 8'h0f, 8'hef, 8'h05, 8'h00, 8'h03, 8'hf1, 8'hfc, 8'h20, 8'h02, 8'hf9, 8'hf4, 8'h19, 8'h03, 8'h01, 8'he4, 8'hf5, 8'h11, 8'hf1, 8'hf5, 8'h06, 8'h0d, 8'hf3, 8'he9, 8'hfa, 8'hed, 8'hec, 8'hed, 8'hf7, 8'hfa, 8'h0c, 8'hfc, 8'h10, 8'hf8, 8'hf4, 8'hdd, 8'hed, 8'hf6, 8'hf9, 8'h01, 8'h18, 8'h16, 8'h04, 8'h1b, 8'h01, 8'h02, 8'hee, 8'hf2, 8'h0c, 8'h0b, 8'h19, 8'hf3, 8'hfb, 8'h15, 8'h17, 8'h0b, 8'he0, 8'h11, 8'h07, 8'hfc, 8'hfb, 8'h14, 8'h09, 8'h17, 8'h05, 8'hea, 8'hf2, 8'he5, 8'he5, 8'h07, 8'hff, 8'h0a, 8'heb, 8'he2, 8'hfa, 8'hfd, 8'h09, 8'h07, 8'h1d},{8'he2, 8'hfd, 8'h00, 8'h04, 8'h11, 8'hec, 8'h10, 8'h0d, 8'hf4, 8'hf7, 8'h17, 8'heb, 8'h13, 8'h00, 8'h0b, 8'h0d, 8'he8, 8'h0f, 8'he1, 8'h01, 8'hff, 8'he7, 8'hfd, 8'h10, 8'hf1, 8'hfa, 8'hfc, 8'h12, 8'h0d, 8'h0a, 8'h03, 8'h04, 8'hdd, 8'hfd, 8'h0b, 8'hf6, 8'hee, 8'h05, 8'h09, 8'hfc, 8'hed, 8'hf6, 8'hf7, 8'hdf, 8'h05, 8'h03, 8'hf0, 8'he7, 8'h15, 8'hef, 8'hff, 8'hf4, 8'hef, 8'h03, 8'h09, 8'h17, 8'hf8, 8'h13, 8'h2d, 8'heb, 8'h10, 8'hfd, 8'h04, 8'h0f, 8'hfc, 8'hf8, 8'h08, 8'h04, 8'h1c, 8'h16, 8'hfd, 8'he4, 8'h18, 8'hf7, 8'h07, 8'hf3, 8'hf9, 8'h10, 8'hed, 8'hf0, 8'h01, 8'h12, 8'hfa, 8'h03, 8'h06, 8'hee, 8'he7, 8'h04, 8'hef, 8'hf7, 8'hfc, 8'he8, 8'h10, 8'h0c, 8'hf6, 8'h04, 8'he6, 8'hf6, 8'he9, 8'hf2, 8'hf3, 8'hfa, 8'he8, 8'h15, 8'h02, 8'h03, 8'he6, 8'h17, 8'heb, 8'h15, 8'h0f, 8'h0c, 8'h16, 8'h00, 8'hdf, 8'hfc, 8'he3, 8'hfe, 8'hfc, 8'hf3, 8'hf9, 8'he5, 8'h0e, 8'hfe, 8'h12, 8'h00, 8'he8, 8'h0d},{8'he3, 8'h0b, 8'he9, 8'h03, 8'hff, 8'hf2, 8'hfa, 8'hec, 8'hf9, 8'hf3, 8'h04, 8'h01, 8'hfa, 8'h1e, 8'h01, 8'h00, 8'hfc, 8'hf5, 8'hf9, 8'h00, 8'hfa, 8'h05, 8'he2, 8'heb, 8'hfb, 8'hf2, 8'hfd, 8'h06, 8'h15, 8'h06, 8'hf8, 8'h13, 8'hee, 8'h12, 8'hff, 8'hfe, 8'he5, 8'h08, 8'h00, 8'hed, 8'h02, 8'he3, 8'h08, 8'hfe, 8'hfd, 8'he0, 8'h18, 8'h02, 8'h01, 8'hf6, 8'h02, 8'h17, 8'h0d, 8'h0a, 8'hec, 8'h11, 8'hf8, 8'hf9, 8'h25, 8'he3, 8'h0e, 8'h16, 8'hf3, 8'hee, 8'hfd, 8'h0e, 8'he5, 8'hf3, 8'h07, 8'h19, 8'hf9, 8'h0d, 8'hf7, 8'hef, 8'h13, 8'hfc, 8'h0a, 8'h12, 8'h02, 8'hf5, 8'h1c, 8'h01, 8'hf8, 8'hf6, 8'h18, 8'h08, 8'h00, 8'h04, 8'h07, 8'h00, 8'h07, 8'he4, 8'h15, 8'he9, 8'hed, 8'h19, 8'hfa, 8'h04, 8'h0b, 8'h13, 8'h17, 8'hec, 8'hfd, 8'hf4, 8'h15, 8'hf2, 8'h0f, 8'h07, 8'he4, 8'hea, 8'hf8, 8'he5, 8'hee, 8'h07, 8'h10, 8'h23, 8'h08, 8'h1e, 8'hea, 8'h02, 8'hed, 8'h0f, 8'h04, 8'hed, 8'hfc, 8'h0a, 8'hfc, 8'h04},{8'hfd, 8'h11, 8'hee, 8'h0c, 8'hea, 8'hee, 8'hf1, 8'hf1, 8'hf7, 8'h0e, 8'h08, 8'h02, 8'hef, 8'he4, 8'h04, 8'hf4, 8'h0d, 8'hf0, 8'h04, 8'hfd, 8'hec, 8'hf7, 8'h07, 8'he5, 8'hfe, 8'hed, 8'h0b, 8'h14, 8'h0f, 8'hfe, 8'hf9, 8'h12, 8'hda, 8'hfc, 8'hee, 8'hf6, 8'hdc, 8'hf5, 8'he7, 8'hf2, 8'hfc, 8'h0a, 8'h1e, 8'hdd, 8'hfa, 8'hfd, 8'h12, 8'h06, 8'h13, 8'h11, 8'hf8, 8'h00, 8'he3, 8'hdf, 8'hf2, 8'h11, 8'he3, 8'hf8, 8'h28, 8'hf3, 8'he9, 8'hfa, 8'hf7, 8'h03, 8'hdf, 8'h06, 8'he8, 8'h0c, 8'h0a, 8'hf5, 8'he7, 8'h07, 8'h15, 8'h0f, 8'hf3, 8'hfd, 8'hf4, 8'hea, 8'hf2, 8'h02, 8'hfe, 8'hf2, 8'he9, 8'h16, 8'hec, 8'he9, 8'h0b, 8'hee, 8'hf0, 8'h07, 8'he1, 8'he4, 8'hec, 8'hf9, 8'hfb, 8'h15, 8'hf2, 8'hf8, 8'h0e, 8'h18, 8'h12, 8'hfb, 8'h16, 8'h09, 8'h10, 8'h00, 8'h0d, 8'h0e, 8'hea, 8'h11, 8'hfb, 8'he2, 8'h01, 8'h00, 8'h05, 8'hec, 8'hf6, 8'hf8, 8'h13, 8'hee, 8'h00, 8'hfb, 8'hdf, 8'h16, 8'hf0, 8'hf8, 8'h18, 8'heb},{8'h0b, 8'h13, 8'h00, 8'h00, 8'he8, 8'h00, 8'h22, 8'h04, 8'hf8, 8'hf0, 8'hf7, 8'hde, 8'heb, 8'hf1, 8'hef, 8'he5, 8'hea, 8'h13, 8'hfc, 8'h1a, 8'h0d, 8'hfd, 8'h07, 8'he5, 8'h06, 8'hd9, 8'hec, 8'hf6, 8'h0b, 8'h16, 8'hde, 8'h18, 8'hef, 8'he8, 8'hf5, 8'h05, 8'hfc, 8'h07, 8'h11, 8'hf1, 8'he9, 8'hee, 8'h10, 8'hf6, 8'h00, 8'h13, 8'h06, 8'h0b, 8'h15, 8'h0a, 8'hff, 8'h10, 8'h14, 8'hfc, 8'hf8, 8'h00, 8'h0f, 8'h04, 8'h21, 8'hf8, 8'hec, 8'hed, 8'hf1, 8'he9, 8'hd8, 8'h06, 8'hdc, 8'hf8, 8'h18, 8'hf4, 8'he5, 8'h0d, 8'h07, 8'h03, 8'h04, 8'h04, 8'hf9, 8'hf0, 8'hfa, 8'h0f, 8'heb, 8'hec, 8'he2, 8'h01, 8'hec, 8'h10, 8'heb, 8'h08, 8'he8, 8'hde, 8'hfe, 8'he5, 8'h1c, 8'h02, 8'h08, 8'h02, 8'h09, 8'he6, 8'he9, 8'hf0, 8'hef, 8'hf3, 8'he7, 8'hfe, 8'hf2, 8'hf0, 8'h17, 8'h0f, 8'he6, 8'hef, 8'hda, 8'hee, 8'hf2, 8'h09, 8'h07, 8'h1e, 8'he3, 8'h04, 8'hec, 8'hdb, 8'h09, 8'h10, 8'hf7, 8'he7, 8'hfe, 8'h03, 8'hee, 8'h0a},};
 assign bias_vector = BIAS_FILE_1;

 always_ff @(posedge clk) begin
        if(rst) begin
    for (k = 0; k < OUT_SIZE_1; k++) 
        output_vector[k] <= '0;
            i <= '0;
        end else begin
            for (k = 0; k < OUT_SIZE_1; k++)
            output_vector[k] <= output_vector_nxt[k];
            i <= i_nxt;
    end
    end
    

    always_comb begin
        
        if (i < IN_SIZE_1) begin
            i_nxt = i + 1;
            for (j = 0; j < OUT_SIZE_1; j++) 
            output_vector_nxt[j] = output_vector[j] +  bias_vector[j] + input_vector[i] * weight_matrix[i][j];
        end else begin
            i_nxt = i;
            for (j = 0; j < OUT_SIZE_1; j++) begin
            if (output_vector[j] < 0) 
            output_vector_nxt [j] = 0;
            else
            output_vector_nxt [j] = output_vector [j];
            end
        end

        end
endmodule
