package ap_parameters;
    //multiplier parameters
    localparam A_WIDTH = 32;
    localparam B_WIDTH = 16;
    localparam P_WIDTH = 32;
    
    endpackage