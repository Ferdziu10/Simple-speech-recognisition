`timescale 1ns / 1ps

module FFT256_tb;

    parameter WIDTH = 16;

    // Testbench signals
    logic                clock;
    logic                reset;
    logic                di_en;
    logic [WIDTH-1:0]    di_re;
    logic [WIDTH-1:0]    di_im;
    logic                do_en;
    logic [WIDTH-1:0]    do_re;
    logic [WIDTH-1:0]    do_im;

    // Instantiate the FFT256 module
    FFT256 #(.WIDTH(WIDTH)) DUT (
        .clock(clock),
        .reset(reset),
        .di_en(di_en),
        .di_re(di_re),
        .di_im(di_im),
        .do_en(do_en),
        .do_re(do_re),
        .do_im(do_im)
    );

    // Clock generation
    always #5 clock = ~clock;

    // Test vectors
    logic [WIDTH-1:0] test_input_re [0:255] = {6314, -5354, -28154, 11432, -24379, 24470, 16680, -15485, -25402, -4122, 31062, -17528, -10346, 4953, -28409, -31515, -31134, 9475, -1484, 30409, -24485, 13112, -26301, 4490, -30570, -21832, -19860, -917, 30846, 13907, -18462, -27496, 28561, -25694, -1342, -8207, 25960, -23490, -22359, 6085, -21681, 8522, -30551, 24961, 15930, 6709, -21999, -5701, 7207, 13753, -3775, -1517, -21149, -21052, 913, 24201, 30281, -19345, -22864, -31014, -18317, -29226, -16530, 13106, 9152, 2293, 29836, 22167, -12912, 29446, 9499, 22840, -16866, 6715, 27506, -20396, -28164, -26554, 1701, 29431, 17609, -30325, 4097, -31176, 23585, -16462, 17290, 11075, 18357, -4017, 14878, -4364, -28302, 8684, 472, 4441, 9304, -32313, -20336, -18326, 25411, -31785, 2472, 18274, 9248, 23536, 4521, 19543, -2258, 8604, 13231, 3584, -5393, 9562, -19916, -14688, -20815, -31689, -24133, -30437, 19274, 1219, -19194, -14888, 21615, 28891, 13034, -22578, 18904, 24447, -24382, -7982, -23392, -4435, -15463, -32261, 22493, -6155, 24579, 16942, -6971, -2880, 2773, 32035, 28631, 6495, -27054, 11326, -2193, -22010, 7861, 6851, -13432, 18016, 29093, -1764, -17931, 15728, 20542, 8723, 27046, 8773, 17977, 6104, 32455, -9757, 20899, -13729, -23303, -13927, 8998, 14874, -27583, -19533, -14080, 25832, 32508, -18589, 26675, -18674, -31631, -30019, -2349, 16015, -5054, 12208, 17917, -30292, 5176, 20471, 8069, -30687, 1222, 16749, -5865, 14632, 23090, 170, 2168, 27302, -29547, 1524, 27999, 3114, -20485, 755, 20957, -11687, 19007, 9107, -11065, -32759, -16018, 12176, -5900, -24508, -6717, 5031, 16972, -22793, -23533, -3079, 8253, 14493, 30074, 12571, 960, 10323, 2951, 9948, -25275, -25441, -30885, -4123, 3651, 28202, -1781, -14890, -22302, -26329, -20743, -24681, -7196, 8743, 2456, 17420, -28056, -31983, 8427, 8637, -23098, -11920, -6577, -2502, 19899, 5589};
    logic [WIDTH-1:0] test_input_im [0:255];
    logic [WIDTH-1:0] expected_output_re [0:255] ={32174, 61611, 62370, 1124, 64718, 3078, 63556, 1493, 3772, 481, 973, 231, 656, 61339, 342, 323, 2601, 64298, 293, 2293, 63501, 62193, 1849, 1027, 2092, 3013, 1860, 2478, 138, 63878, 64224, 58722, 4464, 63551, 62711, 1593, 2950, 760, 1333, 2794, 62683, 1275, 2261, 576, 63345, 2208, 2732, 3384, 2548, 63985, 60262, 63868, 284, 64982, 18, 65232, 64972, 914, 65347, 556, 693, 64382, 513, 65143, 64464, 2405, 2567, 60014, 64323, 63338, 2720, 62628, 3852, 1402, 64429, 64815, 341, 2830, 62951, 64277, 5192, 878, 64591, 64785, 63399, 3035, 64122, 65055, 480, 64535, 65311, 65182, 599, 65174, 2174, 85, 1526, 1860, 2045, 438, 2066, 709, 2211, 62822, 64530, 2580, 1360, 4, 1715, 64555, 63008, 456, 1101, 2765, 62576, 65210, 61883, 63059, 136, 2103, 2960, 64749, 4446, 63966, 64427, 2379, 64066, 62049, 65028, 62049, 64066, 2379, 64427, 63966, 4446, 64749, 2960, 2103, 136, 63059, 61883, 65210, 62576, 2765, 1101, 456, 63008, 64555, 1715, 4, 1360, 2580, 64530, 62822, 2211, 709, 2066, 438, 2045, 1860, 1526, 85, 2174, 65174, 599, 65182, 65311, 64535, 480, 65055, 64122, 3035, 63399, 64785, 64591, 878, 5192, 64277, 62951, 2830, 341, 64815, 64429, 1402, 3852, 62628, 2720, 63338, 64323, 60014, 2567, 2405, 64464, 65143, 513, 64382, 693, 556, 65347, 914, 64972, 65232, 18, 64982, 284, 63868, 60262, 63985, 2548, 3384, 2732, 2208, 63345, 576, 2261, 1275, 62683, 2794, 1333, 760, 2950, 1593, 62711, 63551, 4464, 58722, 64224, 63878, 138, 2478, 1860, 3013, 2092, 1027, 1849, 62193, 63501, 2293, 293, 64298, 2601, 323, 342, 61339, 656, 231, 973, 481, 3772, 1493, 63556, 3078, 64718, 1124, 62370, 61611};
    logic [WIDTH-1:0] expected_output_im [0:255] = {0, 1757, 1056, 700, 63313, 611, 1246, 63083, 62574, 2779, 2474, 2742, 91, 60393, 3678, 60052, 1202, 63943, 942, 64195, 64564, 63435, 2055, 1262, 64169, 64540, 3467, 3960, 1055, 64662, 64370, 452, 139, 63480, 633, 3025, 65335, 883, 64259, 1658, 5630, 1546, 2107, 1682, 439, 1191, 1799, 63714, 2993, 1555, 1853, 4779, 62792, 78, 65399, 4019, 61880, 64820, 63778, 61998, 60517, 4148, 65322, 1013, 64627, 61947, 63231, 2063, 1433, 3141, 65311, 1781, 598, 4944, 1058, 63421, 3471, 3391, 2874, 902, 62266, 1704, 63340, 65455, 65207, 65079, 937, 282, 201, 63903, 1006, 63162, 64844, 1141, 63087, 389, 65476, 1441, 63656, 2982, 63479, 62183, 64095, 2100, 64693, 64348, 65192, 64809, 61552, 2210, 64259, 62414, 64760, 63395, 63891, 365, 62512, 3263, 4606, 65425, 64420, 65527, 814, 63609, 65436, 64909, 63844, 222, 0, 65314, 1692, 627, 100, 1927, 64722, 9, 1116, 111, 60930, 62273, 3024, 65171, 1645, 2141, 776, 3122, 1277, 63326, 3984, 727, 344, 1188, 843, 63436, 1441, 3353, 2057, 62554, 1880, 64095, 60, 65147, 2449, 64395, 692, 2374, 64530, 1633, 65335, 65254, 64599, 457, 329, 81, 2196, 63832, 3270, 64634, 62662, 62145, 62065, 2115, 64478, 60592, 64938, 63755, 225, 62395, 64103, 63473, 2305, 3589, 909, 64523, 214, 61388, 5019, 3538, 1758, 716, 3656, 61517, 137, 65458, 2744, 60757, 63683, 63981, 62543, 1822, 63737, 64345, 65097, 63854, 63429, 63990, 59906, 63878, 1277, 64653, 201, 62511, 64903, 2056, 65397, 65084, 1166, 874, 64481, 61576, 62069, 996, 1367, 64274, 63481, 2101, 972, 1341, 64594, 1593, 64334, 5484, 61858, 5143, 65445, 62794, 63062, 62757, 2962, 2453, 64290, 64925, 2223, 64836, 64480, 63779};

    integer i;

    initial begin
        for (i = 0; i < 256; i = i + 1) 
            test_input_im[i] = 0;
        // Initialize signals
        clock = 0;
        reset = 1;
        di_en = 0;
        di_re = 0;
        di_im = 0;

  

        // Release reset
        #15 reset = 0;

        // Apply input data
        for (i = 0; i < 256; i = i + 1) begin
            #10;
            di_en = 1;
            di_re = test_input_re[i];
            di_im = test_input_im[i];
        end
        di_en = 0;


        // Wait for FFT output
        #50000;

        // Check output data
        for (i = 0; i < 256; i = i + 1) begin
            #10;
            if (do_en) begin
                if (do_re !== expected_output_re[i] || do_im !== expected_output_im[i]) begin
                    $display("ERROR: Output mismatch at index %d: Expected (%d, %d), Got (%d, %d)",
                        i, expected_output_re[i], expected_output_im[i], do_re, do_im);
                end else begin
                    $display("PASS: Output match at index %d: (%d, %d)",
                        i, do_re, do_im);
                end
            end
        end

        // End simulation
        $finish;
    end
endmodule