import nn_parameters::*;

module dense_layer_2 (
    input clk,
    input rst,
    input logic signed [23:0] input_vector [IN_SIZE_2-1:0],
    output logic signed [31:0] output_vector [OUT_SIZE_2-1:0]
);


    logic signed [7:0] weight_matrix [IN_SIZE_2-1:0][OUT_SIZE_2-1:0];
    logic signed [7:0] bias_vector [OUT_SIZE_2-1:0];
    logic signed [31:0] output_vector_nxt [OUT_SIZE_2-1:0];
    logic [7:0] i;
    logic [7:0] i_nxt;

    integer j, k;

assign weight_matrix[0] = {8'hed, 8'hf9, 8'h06, 8'hf6, 8'hf6, 8'hf9, 8'h0a, 8'hf9, 8'hf8, 8'h14, 8'h0a, 8'h04, 8'hfb, 8'h00, 8'h0b, 8'h05, 8'h13, 8'hea, 8'hf3, 8'h12, 8'h07, 8'hfb, 8'h01, 8'h13, 8'h0a, 8'h03, 8'h11, 8'hfa, 8'h03, 8'h10, 8'hf1, 8'h00, 8'h10, 8'hf5, 8'hf7, 8'hf3, 8'h10, 8'he7, 8'hff, 8'h02, 8'he9, 8'hf8, 8'h0c, 8'h04, 8'he6, 8'hea, 8'h11, 8'hf3, 8'hf1, 8'hf9, 8'h02, 8'h05, 8'h0f, 8'hfd, 8'h06, 8'h07, 8'hfb, 8'h01, 8'he3, 8'h13, 8'hf4, 8'hf1, 8'hfe, 8'h0d};
assign weight_matrix[1] = {8'h00, 8'hf7, 8'hf1, 8'hf4, 8'hf8, 8'h02, 8'h05, 8'hf5, 8'hfe, 8'h05, 8'hf2, 8'hf0, 8'hff, 8'h16, 8'hfb, 8'h04, 8'h0f, 8'h06, 8'h05, 8'h05, 8'hea, 8'h12, 8'h0d, 8'h01, 8'h06, 8'h10, 8'hff, 8'hec, 8'hfb, 8'hfc, 8'h09, 8'h06, 8'h07, 8'hfb, 8'hfa, 8'h06, 8'hf6, 8'h13, 8'hf1, 8'hef, 8'h15, 8'hf7, 8'h05, 8'h08, 8'hfc, 8'hf8, 8'h15, 8'hec, 8'hfa, 8'hf0, 8'hf6, 8'hfc, 8'hfa, 8'hf5, 8'h10, 8'hed, 8'h13, 8'hff, 8'h15, 8'hfc, 8'hfb, 8'hf3, 8'hfb, 8'h0b};
assign weight_matrix[2] = {8'h01, 8'hf2, 8'h04, 8'hee, 8'h03, 8'h02, 8'hf6, 8'hf3, 8'h00, 8'h0e, 8'h0b, 8'hf9, 8'h0a, 8'hf7, 8'h10, 8'h0b, 8'hf2, 8'hff, 8'hfa, 8'hf2, 8'heb, 8'hfe, 8'hf0, 8'hed, 8'he8, 8'h02, 8'hee, 8'h0f, 8'hf0, 8'heb, 8'h10, 8'h09, 8'hfc, 8'h0b, 8'h0a, 8'hf6, 8'h04, 8'h05, 8'h14, 8'hf7, 8'he9, 8'h07, 8'h0c, 8'h0d, 8'h00, 8'hfd, 8'hec, 8'hf7, 8'hf4, 8'hfc, 8'h0a, 8'hf3, 8'hf9, 8'h07, 8'hf7, 8'h0a, 8'h14, 8'h09, 8'h03, 8'h0a, 8'he9, 8'h0e, 8'h02, 8'hfd};
assign weight_matrix[3] = {8'hfa, 8'h14, 8'hf5, 8'he7, 8'hea, 8'h0e, 8'h20, 8'h10, 8'h0d, 8'hf1, 8'hf2, 8'h04, 8'hf3, 8'hf0, 8'hf5, 8'heb, 8'hf9, 8'hfb, 8'h08, 8'h00, 8'h09, 8'h09, 8'he9, 8'h0c, 8'h0d, 8'h06, 8'he9, 8'h0c, 8'hfd, 8'hef, 8'hf4, 8'h09, 8'heb, 8'h0c, 8'h06, 8'h12, 8'hf3, 8'h10, 8'hfe, 8'hf1, 8'hee, 8'hf5, 8'hfa, 8'hf5, 8'h12, 8'h0f, 8'hf0, 8'hf8, 8'hec, 8'hed, 8'h09, 8'h00, 8'h01, 8'he7, 8'h02, 8'he9, 8'hfb, 8'hfc, 8'hec, 8'hfc, 8'hf3, 8'hff, 8'h05, 8'h02};
assign weight_matrix[4] = {8'h05, 8'h14, 8'he2, 8'hfb, 8'h03, 8'he4, 8'h04, 8'h06, 8'hf9, 8'hfe, 8'hf6, 8'h08, 8'h07, 8'hfb, 8'he8, 8'heb, 8'h0c, 8'hf5, 8'h13, 8'hed, 8'h11, 8'h08, 8'hef, 8'hed, 8'h07, 8'h0a, 8'h09, 8'he9, 8'h07, 8'hf9, 8'he4, 8'h12, 8'hf4, 8'h04, 8'he8, 8'hf5, 8'he6, 8'h09, 8'hf6, 8'hf6, 8'hf7, 8'h11, 8'hef, 8'h15, 8'hf7, 8'hfe, 8'h06, 8'h04, 8'hf3, 8'he7, 8'hfe, 8'h19, 8'hee, 8'hfd, 8'hf7, 8'he3, 8'hf5, 8'hf9, 8'h04, 8'hf2, 8'h0e, 8'hfe, 8'h16, 8'hf0};
assign weight_matrix[5] = {8'hf1, 8'h0d, 8'h02, 8'hfc, 8'hf0, 8'hfb, 8'hf6, 8'h13, 8'hee, 8'hed, 8'hf1, 8'h07, 8'hfe, 8'hf5, 8'h11, 8'h02, 8'h0c, 8'h08, 8'h03, 8'h12, 8'hf7, 8'h09, 8'hf1, 8'hf9, 8'h01, 8'h1c, 8'h06, 8'h08, 8'h13, 8'h07, 8'hf3, 8'h11, 8'hf4, 8'hf9, 8'h10, 8'hea, 8'hec, 8'hf5, 8'h13, 8'h10, 8'h04, 8'hfd, 8'hef, 8'h11, 8'h0d, 8'hfd, 8'h00, 8'h0b, 8'h0f, 8'hee, 8'hf7, 8'h0d, 8'h0a, 8'hf9, 8'hf7, 8'h0d, 8'h09, 8'h00, 8'h10, 8'hfe, 8'h05, 8'h0c, 8'hf8, 8'hfe};
assign weight_matrix[6] = {8'he8, 8'h12, 8'h0f, 8'hfa, 8'hf6, 8'hfc, 8'he5, 8'h05, 8'hf0, 8'hf3, 8'hfd, 8'hf2, 8'h03, 8'h0c, 8'hff, 8'hff, 8'h14, 8'hee, 8'h00, 8'h0a, 8'h08, 8'hfd, 8'h05, 8'hed, 8'hf7, 8'hf8, 8'he8, 8'h0f, 8'h11, 8'h00, 8'he8, 8'h03, 8'h10, 8'h0c, 8'h08, 8'h06, 8'hfb, 8'hf1, 8'he9, 8'h06, 8'hfc, 8'h0f, 8'hf9, 8'hf5, 8'hf3, 8'h13, 8'hfe, 8'hff, 8'h12, 8'h10, 8'h0d, 8'hed, 8'h12, 8'hf6, 8'h08, 8'hf8, 8'hf6, 8'h20, 8'h0a, 8'hee, 8'hfa, 8'h1a, 8'hf3, 8'h04};
assign weight_matrix[7] = {8'h04, 8'hea, 8'h09, 8'h05, 8'hf0, 8'hec, 8'hfd, 8'h07, 8'hfe, 8'hf2, 8'h14, 8'h12, 8'h0e, 8'hfb, 8'h02, 8'h0f, 8'h0d, 8'h0d, 8'heb, 8'h07, 8'h04, 8'hec, 8'h01, 8'hf4, 8'h09, 8'hfa, 8'hf5, 8'h00, 8'hf3, 8'hf8, 8'h12, 8'hf4, 8'heb, 8'h08, 8'hf5, 8'hfd, 8'hf4, 8'hf2, 8'hf0, 8'hf3, 8'h12, 8'hf5, 8'h0c, 8'hf5, 8'hed, 8'h13, 8'hef, 8'he7, 8'h13, 8'hf5, 8'hf8, 8'h03, 8'h04, 8'hf8, 8'heb, 8'hf9, 8'hee, 8'hf1, 8'h14, 8'h07, 8'h05, 8'h07, 8'h02, 8'h13};
assign weight_matrix[8] = {8'hf5, 8'he4, 8'h0e, 8'hf4, 8'h13, 8'hfa, 8'hf2, 8'hf1, 8'hfb, 8'hed, 8'hff, 8'hf9, 8'hf4, 8'hfd, 8'h02, 8'h0a, 8'hfa, 8'h00, 8'h0a, 8'h02, 8'hef, 8'hfe, 8'hfd, 8'h0c, 8'he7, 8'hd7, 8'h06, 8'hfa, 8'hf5, 8'hfd, 8'hfd, 8'hf4, 8'h11, 8'h02, 8'h12, 8'hf8, 8'hf9, 8'hfe, 8'he7, 8'h0a, 8'h0a, 8'h1a, 8'h0b, 8'h05, 8'h06, 8'h0b, 8'hf4, 8'hfb, 8'h01, 8'hef, 8'h13, 8'hfd, 8'hf2, 8'heb, 8'h12, 8'h07, 8'hfa, 8'hf7, 8'he7, 8'h0f, 8'h07, 8'he7, 8'hfa, 8'h07};
assign weight_matrix[9] = {8'hfc, 8'h10, 8'h0f, 8'hed, 8'h14, 8'hed, 8'h11, 8'hed, 8'h13, 8'h0e, 8'hf6, 8'hf5, 8'h07, 8'h00, 8'hf4, 8'h0c, 8'h08, 8'hf8, 8'hea, 8'h02, 8'h16, 8'h10, 8'h0f, 8'h14, 8'hfe, 8'hf7, 8'hf4, 8'hf2, 8'hf7, 8'h16, 8'h06, 8'hff, 8'h0f, 8'hea, 8'h15, 8'hff, 8'h13, 8'hff, 8'h07, 8'hfa, 8'hef, 8'h00, 8'hef, 8'hf5, 8'h12, 8'hf3, 8'h0e, 8'heb, 8'hfe, 8'h06, 8'hef, 8'h07, 8'hed, 8'hf4, 8'hee, 8'hea, 8'h03, 8'h0e, 8'hf3, 8'hec, 8'h01, 8'hf4, 8'h12, 8'h0c};
assign weight_matrix[10] = {8'h04, 8'hef, 8'hfa, 8'hff, 8'h09, 8'h07, 8'hf0, 8'hf9, 8'hf9, 8'hf1, 8'hff, 8'h09, 8'hfd, 8'hf5, 8'h16, 8'h02, 8'hf4, 8'h0b, 8'hec, 8'h08, 8'hf8, 8'h09, 8'h02, 8'hef, 8'h00, 8'h01, 8'h06, 8'h12, 8'h0c, 8'h11, 8'hea, 8'h13, 8'heb, 8'hff, 8'h14, 8'h09, 8'hf7, 8'h15, 8'h13, 8'h15, 8'h04, 8'h15, 8'h02, 8'h05, 8'h15, 8'hfa, 8'h0c, 8'h12, 8'hf9, 8'hf8, 8'h0a, 8'h03, 8'h09, 8'h01, 8'hf7, 8'h12, 8'h05, 8'hf0, 8'h07, 8'h0c, 8'hfb, 8'h0d, 8'h11, 8'h0a};
assign weight_matrix[11] = {8'h0f, 8'h0c, 8'h0f, 8'hed, 8'hf1, 8'he8, 8'hec, 8'hf2, 8'hfb, 8'h06, 8'hf5, 8'hf5, 8'h06, 8'h0a, 8'h10, 8'h10, 8'hea, 8'hf2, 8'hfa, 8'h03, 8'h02, 8'h06, 8'hff, 8'h11, 8'h05, 8'h06, 8'h12, 8'hf7, 8'h05, 8'h05, 8'hec, 8'h11, 8'h01, 8'h03, 8'h11, 8'h02, 8'h10, 8'h07, 8'h0b, 8'hec, 8'h00, 8'hfc, 8'hff, 8'h0b, 8'hf7, 8'h02, 8'h0a, 8'h12, 8'hec, 8'hf7, 8'h09, 8'h12, 8'hfc, 8'hfa, 8'heb, 8'h10, 8'h0d, 8'h02, 8'h02, 8'hfb, 8'h12, 8'h12, 8'h08, 8'hf5};
assign weight_matrix[12] = {8'h11, 8'hf9, 8'heb, 8'h00, 8'h09, 8'h00, 8'h1d, 8'hef, 8'hf7, 8'hed, 8'hfa, 8'hf2, 8'h16, 8'hf7, 8'h12, 8'hfe, 8'hff, 8'h10, 8'h20, 8'hef, 8'h0b, 8'hf2, 8'hfb, 8'hfb, 8'h05, 8'hd4, 8'hfb, 8'hfd, 8'hf9, 8'hef, 8'h08, 8'h1a, 8'hdf, 8'h00, 8'hf0, 8'hf4, 8'h0b, 8'hef, 8'h0f, 8'h02, 8'he6, 8'hea, 8'hf2, 8'h15, 8'h04, 8'h13, 8'hf6, 8'hf3, 8'hfa, 8'h0c, 8'he7, 8'h10, 8'h10, 8'hfb, 8'he1, 8'hff, 8'hfd, 8'hde, 8'hf5, 8'hfc, 8'hf7, 8'he8, 8'h24, 8'h36};
assign weight_matrix[13] = {8'h08, 8'h01, 8'h07, 8'h0c, 8'hf1, 8'h05, 8'hf5, 8'hf2, 8'h0c, 8'hfa, 8'hf0, 8'h0f, 8'hf2, 8'hef, 8'hfe, 8'h0a, 8'hf6, 8'hf5, 8'h02, 8'h02, 8'hfb, 8'h14, 8'h06, 8'hf8, 8'h0e, 8'h0f, 8'h12, 8'hec, 8'heb, 8'h09, 8'h0c, 8'hf6, 8'h0d, 8'hf0, 8'hfc, 8'hed, 8'h09, 8'he8, 8'hfa, 8'h0a, 8'hf9, 8'h0c, 8'hff, 8'hfc, 8'he9, 8'hf4, 8'h08, 8'h11, 8'hf8, 8'hf2, 8'hf9, 8'hef, 8'h01, 8'hfb, 8'h0f, 8'hfa, 8'hf6, 8'hf7, 8'hf2, 8'h0f, 8'h06, 8'h11, 8'h00, 8'he9};
assign weight_matrix[14] = {8'hec, 8'h16, 8'hfc, 8'hff, 8'h13, 8'h0d, 8'hf0, 8'hf3, 8'hfd, 8'hfe, 8'h13, 8'hf8, 8'hec, 8'hf2, 8'hed, 8'h0c, 8'h03, 8'h00, 8'h05, 8'hfe, 8'hef, 8'h06, 8'hea, 8'h06, 8'hf6, 8'h00, 8'hfd, 8'h06, 8'h11, 8'hec, 8'h0f, 8'h10, 8'h10, 8'h0b, 8'hf7, 8'hf2, 8'h02, 8'h15, 8'h13, 8'hec, 8'hf8, 8'hf0, 8'hf4, 8'hfa, 8'hff, 8'hec, 8'h0f, 8'h16, 8'hf4, 8'hf9, 8'h04, 8'h04, 8'hed, 8'h0a, 8'h12, 8'hed, 8'h08, 8'h12, 8'hf7, 8'h06, 8'hf7, 8'hf3, 8'h0a, 8'h10};
assign weight_matrix[15] = {8'h03, 8'h0a, 8'hf9, 8'h17, 8'h13, 8'h0c, 8'hfb, 8'h01, 8'h08, 8'hed, 8'hf9, 8'h08, 8'hf5, 8'hfd, 8'h09, 8'h10, 8'hf0, 8'h06, 8'h06, 8'hf1, 8'h02, 8'hff, 8'hf5, 8'he2, 8'hed, 8'h02, 8'h04, 8'h10, 8'heb, 8'hf4, 8'h09, 8'h1d, 8'hd6, 8'h08, 8'h10, 8'h11, 8'h1e, 8'h1c, 8'h0a, 8'hfc, 8'hf6, 8'h02, 8'hec, 8'hfb, 8'h03, 8'h17, 8'h03, 8'he9, 8'hdf, 8'he8, 8'hfc, 8'h16, 8'hf4, 8'h27, 8'h04, 8'heb, 8'h03, 8'hef, 8'hf7, 8'hee, 8'h01, 8'h00, 8'h0c, 8'h00};
assign weight_matrix[16] = {8'h02, 8'hea, 8'h11, 8'hee, 8'h11, 8'h12, 8'hf8, 8'h07, 8'h01, 8'h16, 8'h14, 8'hef, 8'h08, 8'h02, 8'h0e, 8'hfb, 8'hfb, 8'hf0, 8'hf7, 8'hec, 8'hf1, 8'hf9, 8'hfa, 8'hf0, 8'hfa, 8'h0c, 8'h12, 8'hf6, 8'h08, 8'h05, 8'h03, 8'hf9, 8'hf3, 8'h0b, 8'heb, 8'heb, 8'hec, 8'hfe, 8'h01, 8'heb, 8'hec, 8'hf3, 8'hf2, 8'hf2, 8'hfc, 8'h09, 8'h04, 8'h03, 8'hfc, 8'h0b, 8'hee, 8'hfc, 8'h16, 8'hf7, 8'h03, 8'hfd, 8'h04, 8'h11, 8'h15, 8'h0d, 8'h16, 8'hf1, 8'h0e, 8'hec};
assign weight_matrix[17] = {8'h10, 8'hfd, 8'hfa, 8'hfe, 8'hfb, 8'hee, 8'hfb, 8'hf6, 8'h0d, 8'h0b, 8'h13, 8'h14, 8'hf2, 8'h04, 8'hfa, 8'h03, 8'h07, 8'h01, 8'h04, 8'hef, 8'h0b, 8'hf4, 8'h00, 8'h15, 8'hf9, 8'hec, 8'h05, 8'hf7, 8'h12, 8'hf3, 8'hec, 8'h11, 8'h11, 8'h0d, 8'hfe, 8'hf4, 8'hfc, 8'h11, 8'hec, 8'h0e, 8'h0b, 8'hea, 8'hf4, 8'hff, 8'h04, 8'hea, 8'hec, 8'hfe, 8'h00, 8'h08, 8'hea, 8'hfe, 8'hf7, 8'h12, 8'hf6, 8'hfc, 8'hef, 8'h0b, 8'hf5, 8'hed, 8'h0f, 8'hf6, 8'hf9, 8'hfb};
assign weight_matrix[18] = {8'heb, 8'hef, 8'hfb, 8'hf7, 8'hf5, 8'hec, 8'h07, 8'hee, 8'hfa, 8'hf7, 8'hf6, 8'h05, 8'h11, 8'h0f, 8'hfd, 8'hfb, 8'hf7, 8'hf9, 8'h12, 8'h10, 8'hee, 8'h0c, 8'hf5, 8'hed, 8'h0c, 8'hfa, 8'he8, 8'hf6, 8'hfc, 8'h08, 8'h02, 8'hed, 8'hfc, 8'h0c, 8'hee, 8'h04, 8'hee, 8'hf8, 8'hf6, 8'he9, 8'hfd, 8'hed, 8'h05, 8'hf5, 8'hf8, 8'h10, 8'hfa, 8'hf6, 8'hfb, 8'hef, 8'hf3, 8'h0e, 8'h0e, 8'hec, 8'hf2, 8'h0c, 8'hfb, 8'h02, 8'hf8, 8'hf3, 8'hf3, 8'hfb, 8'hf5, 8'h0b};
assign weight_matrix[19] = {8'h06, 8'hf2, 8'h0d, 8'he7, 8'hfb, 8'hf0, 8'h13, 8'hec, 8'hf3, 8'h0c, 8'hef, 8'h08, 8'h08, 8'h00, 8'hf4, 8'hfc, 8'h12, 8'hf0, 8'hfb, 8'hfc, 8'h02, 8'h04, 8'hf1, 8'h01, 8'he9, 8'h08, 8'hee, 8'hf0, 8'hf2, 8'h11, 8'hff, 8'heb, 8'hf6, 8'hf3, 8'h0b, 8'h09, 8'h09, 8'h0b, 8'hf0, 8'h05, 8'hf5, 8'hfc, 8'h0c, 8'h00, 8'hf6, 8'h02, 8'hf9, 8'h04, 8'h0a, 8'hff, 8'h12, 8'hfa, 8'hf8, 8'h04, 8'hf4, 8'hed, 8'hef, 8'h0f, 8'hf5, 8'h08, 8'hf2, 8'h08, 8'hf6, 8'h0b};
assign weight_matrix[20] = {8'h13, 8'hf9, 8'hf0, 8'h10, 8'hed, 8'hf5, 8'h12, 8'hf6, 8'h00, 8'h07, 8'hea, 8'heb, 8'h10, 8'h14, 8'h13, 8'h10, 8'hf0, 8'hf0, 8'hfe, 8'h05, 8'h0f, 8'h10, 8'hf7, 8'hf7, 8'hef, 8'h11, 8'h04, 8'hf1, 8'h09, 8'h12, 8'h02, 8'h01, 8'hf9, 8'h13, 8'hfc, 8'h09, 8'hee, 8'h09, 8'h11, 8'h0e, 8'h06, 8'h11, 8'h0f, 8'h13, 8'h0e, 8'hf1, 8'hf1, 8'h12, 8'hf2, 8'h0b, 8'h02, 8'hf6, 8'h0a, 8'hee, 8'h0a, 8'h0e, 8'h00, 8'hf5, 8'h0e, 8'hfb, 8'h16, 8'h11, 8'hf7, 8'hf3};
assign weight_matrix[21] = {8'h16, 8'h05, 8'h0a, 8'hfe, 8'hfb, 8'hf8, 8'hf6, 8'hf9, 8'h09, 8'hfb, 8'h0d, 8'hfe, 8'h06, 8'hf4, 8'hff, 8'h08, 8'hfa, 8'hf1, 8'hf7, 8'h0a, 8'h16, 8'h16, 8'hfb, 8'hf1, 8'hf6, 8'hee, 8'h09, 8'hfe, 8'hf7, 8'hfa, 8'h04, 8'hec, 8'hfe, 8'hf4, 8'hee, 8'h11, 8'hff, 8'h06, 8'hf7, 8'hf5, 8'h0c, 8'h16, 8'h02, 8'h0c, 8'h0b, 8'h04, 8'hf5, 8'hfb, 8'h14, 8'h0b, 8'hf5, 8'h15, 8'hfd, 8'h11, 8'h05, 8'h0b, 8'h02, 8'heb, 8'h14, 8'h14, 8'hed, 8'h09, 8'h16, 8'h0f};
assign weight_matrix[22] = {8'h03, 8'heb, 8'h0e, 8'h11, 8'hf7, 8'h06, 8'h01, 8'heb, 8'h04, 8'h0c, 8'hf4, 8'h08, 8'hfc, 8'hf9, 8'h10, 8'h06, 8'h11, 8'h05, 8'hf3, 8'h13, 8'hf6, 8'hf3, 8'h11, 8'h08, 8'h0b, 8'hf2, 8'h0a, 8'hfd, 8'h01, 8'h07, 8'hfb, 8'hf1, 8'hee, 8'hfc, 8'h0c, 8'hfb, 8'h0b, 8'hf6, 8'h0e, 8'h10, 8'he7, 8'hfa, 8'hf3, 8'hf8, 8'h11, 8'hf5, 8'hf6, 8'h0e, 8'h0c, 8'h11, 8'hf0, 8'hef, 8'h00, 8'hef, 8'hf5, 8'h0a, 8'h01, 8'h0c, 8'heb, 8'h08, 8'hf8, 8'hf6, 8'h0c, 8'hfd};
assign weight_matrix[23] = {8'h0d, 8'hfc, 8'hee, 8'h0c, 8'hee, 8'hfc, 8'hfe, 8'h10, 8'h14, 8'he9, 8'h00, 8'he9, 8'h0a, 8'hf8, 8'h05, 8'h0c, 8'h10, 8'h06, 8'h06, 8'h06, 8'hf4, 8'h03, 8'h0c, 8'h08, 8'hf4, 8'hfd, 8'hfc, 8'hf0, 8'hea, 8'h12, 8'heb, 8'h0e, 8'h0f, 8'h06, 8'he8, 8'h14, 8'h0f, 8'hf3, 8'h08, 8'hf9, 8'hf9, 8'hf6, 8'hf3, 8'h0f, 8'h05, 8'hf9, 8'h04, 8'h01, 8'hef, 8'hf6, 8'h0e, 8'h11, 8'hfc, 8'hea, 8'hf4, 8'h01, 8'h0f, 8'h0d, 8'hef, 8'hf9, 8'hf6, 8'hef, 8'h0a, 8'h03};
assign weight_matrix[24] = {8'h0b, 8'hf6, 8'hf0, 8'hf2, 8'h06, 8'h02, 8'h05, 8'h14, 8'hff, 8'hea, 8'h10, 8'h12, 8'hef, 8'h12, 8'h10, 8'h13, 8'hf4, 8'hfb, 8'hfb, 8'h0d, 8'hfd, 8'h15, 8'h14, 8'h0f, 8'hec, 8'h02, 8'h06, 8'hf5, 8'h10, 8'h14, 8'h06, 8'h08, 8'hf4, 8'hff, 8'h0a, 8'hee, 8'h0f, 8'h14, 8'h16, 8'hf5, 8'hf8, 8'hf7, 8'heb, 8'h0f, 8'h0d, 8'hfc, 8'hf4, 8'hfb, 8'hf4, 8'hf6, 8'hec, 8'hfb, 8'h0d, 8'h14, 8'h0a, 8'hfd, 8'h03, 8'h0e, 8'hf4, 8'hea, 8'hf5, 8'h09, 8'hfc, 8'h05};
assign weight_matrix[25] = {8'h0c, 8'he6, 8'hf0, 8'h07, 8'h04, 8'hff, 8'h2e, 8'hfe, 8'hf5, 8'hdf, 8'heb, 8'h05, 8'h1b, 8'he5, 8'hf5, 8'hf8, 8'hff, 8'hf4, 8'h24, 8'hf8, 8'h00, 8'hf4, 8'hfb, 8'hde, 8'hf3, 8'hf9, 8'h04, 8'h10, 8'hed, 8'hd2, 8'hf7, 8'h39, 8'hf8, 8'hfc, 8'h03, 8'hef, 8'hfe, 8'h0b, 8'h18, 8'hf0, 8'hef, 8'h15, 8'hf5, 8'h1a, 8'hea, 8'h0c, 8'hff, 8'h05, 8'h0b, 8'h14, 8'hee, 8'h2b, 8'hf9, 8'hff, 8'hfb, 8'h09, 8'he4, 8'he7, 8'hfd, 8'h0c, 8'h09, 8'hfc, 8'h17, 8'h15};
assign weight_matrix[26] = {8'h06, 8'h11, 8'h0d, 8'h16, 8'hfb, 8'hfc, 8'h09, 8'h10, 8'h0b, 8'hf8, 8'h0f, 8'hf6, 8'h00, 8'hf6, 8'hfc, 8'h11, 8'hf2, 8'h10, 8'h0e, 8'h14, 8'h13, 8'hfb, 8'h12, 8'h12, 8'hec, 8'hed, 8'h0b, 8'hea, 8'h11, 8'h0f, 8'h0b, 8'h07, 8'heb, 8'h07, 8'h13, 8'h0f, 8'h02, 8'h08, 8'h04, 8'h09, 8'h09, 8'h12, 8'h0f, 8'hff, 8'h10, 8'h05, 8'hf5, 8'hf0, 8'hed, 8'h01, 8'h16, 8'h00, 8'h09, 8'h14, 8'h09, 8'h0a, 8'h0f, 8'hff, 8'hf4, 8'hf7, 8'hfe, 8'h05, 8'h0f, 8'hff};
assign weight_matrix[27] = {8'h03, 8'hec, 8'hf9, 8'hf6, 8'h15, 8'h0c, 8'hf0, 8'h14, 8'hec, 8'hf4, 8'h13, 8'h03, 8'h0b, 8'hef, 8'hfd, 8'he9, 8'hec, 8'h0c, 8'hee, 8'hfb, 8'h0b, 8'h06, 8'hf3, 8'h05, 8'hed, 8'hf3, 8'h0f, 8'heb, 8'h0c, 8'h14, 8'h0f, 8'hf4, 8'h0b, 8'heb, 8'h10, 8'h13, 8'hfd, 8'hee, 8'h02, 8'h06, 8'h08, 8'h11, 8'h02, 8'hef, 8'h12, 8'hf1, 8'hf6, 8'hf8, 8'hff, 8'hf6, 8'hed, 8'h0f, 8'h00, 8'h08, 8'h14, 8'h14, 8'hff, 8'h04, 8'h0c, 8'hf8, 8'hfc, 8'h10, 8'h00, 8'h02};
assign weight_matrix[28] = {8'hef, 8'h15, 8'h00, 8'he7, 8'h10, 8'h09, 8'hfc, 8'hf5, 8'h01, 8'hf9, 8'h0d, 8'h01, 8'h05, 8'h09, 8'h05, 8'h0a, 8'h04, 8'hf8, 8'h02, 8'h0c, 8'hf4, 8'h0b, 8'h12, 8'hf4, 8'h00, 8'h03, 8'heb, 8'hfb, 8'h01, 8'h02, 8'h0d, 8'hf5, 8'h01, 8'hf8, 8'hea, 8'h13, 8'hfd, 8'hf5, 8'h00, 8'hfc, 8'hef, 8'hff, 8'h0f, 8'hf2, 8'he9, 8'h04, 8'hee, 8'h07, 8'h05, 8'hee, 8'h0a, 8'h02, 8'hf3, 8'hf7, 8'h13, 8'h11, 8'hfb, 8'hff, 8'hf8, 8'hea, 8'h0c, 8'h0d, 8'hf6, 8'hf0};
assign weight_matrix[29] = {8'h05, 8'he8, 8'h10, 8'hee, 8'hf5, 8'hf7, 8'h06, 8'hf1, 8'h1a, 8'h05, 8'hf9, 8'h0a, 8'h10, 8'he8, 8'h1b, 8'h1a, 8'hff, 8'he6, 8'h14, 8'hf6, 8'h0b, 8'hfe, 8'h14, 8'he8, 8'h0c, 8'h0f, 8'h16, 8'hf5, 8'hfd, 8'hec, 8'h05, 8'h26, 8'h08, 8'hf8, 8'hec, 8'hed, 8'h17, 8'hf9, 8'hee, 8'he7, 8'hf6, 8'hfe, 8'h05, 8'h25, 8'h10, 8'h11, 8'hfd, 8'hec, 8'h11, 8'h08, 8'hf0, 8'hf4, 8'h02, 8'h01, 8'hf8, 8'hed, 8'h0a, 8'hf7, 8'hf9, 8'h11, 8'h17, 8'hdf, 8'h22, 8'h2b};
assign weight_matrix[30] = {8'h03, 8'hf5, 8'hf9, 8'h0b, 8'hfb, 8'hf4, 8'hf9, 8'hf4, 8'h03, 8'hf4, 8'h04, 8'h13, 8'h16, 8'hea, 8'h01, 8'he9, 8'hff, 8'hed, 8'hfa, 8'he6, 8'hfa, 8'h03, 8'hf8, 8'hf8, 8'hf5, 8'hd6, 8'hf0, 8'he3, 8'hf9, 8'hfc, 8'h09, 8'h00, 8'hf7, 8'hfe, 8'hf6, 8'hed, 8'he3, 8'he9, 8'hf6, 8'h07, 8'hf1, 8'hf4, 8'hf2, 8'h02, 8'hf2, 8'hfe, 8'hf8, 8'h07, 8'he4, 8'hec, 8'hf5, 8'hfc, 8'h05, 8'hea, 8'h03, 8'hea, 8'hed, 8'hd6, 8'hf9, 8'hfd, 8'h02, 8'he4, 8'h15, 8'h13};
assign weight_matrix[31] = {8'hfe, 8'hf8, 8'h15, 8'hf7, 8'hfd, 8'heb, 8'h0c, 8'hf7, 8'h02, 8'h15, 8'hfd, 8'hfc, 8'hf6, 8'h15, 8'h0e, 8'hf7, 8'hee, 8'h11, 8'h0e, 8'hfd, 8'h0b, 8'hf9, 8'h07, 8'hfc, 8'h14, 8'hed, 8'hfb, 8'hf7, 8'hff, 8'hf2, 8'h05, 8'hf8, 8'h0b, 8'hf3, 8'h14, 8'h07, 8'h15, 8'h12, 8'h16, 8'h16, 8'hfe, 8'h06, 8'h0e, 8'hfb, 8'h0e, 8'h0f, 8'hea, 8'hea, 8'h11, 8'hf8, 8'h14, 8'h00, 8'heb, 8'hf6, 8'h16, 8'h00, 8'hfa, 8'hf2, 8'h16, 8'h16, 8'h01, 8'hf4, 8'hec, 8'hfc};
assign weight_matrix[32] = {8'h0a, 8'hfa, 8'he9, 8'hff, 8'h01, 8'h0c, 8'hfc, 8'h0b, 8'heb, 8'h0c, 8'h14, 8'h03, 8'hfe, 8'h0a, 8'h06, 8'h0e, 8'hed, 8'hf1, 8'h01, 8'hfd, 8'h12, 8'heb, 8'hf3, 8'h06, 8'h0b, 8'h03, 8'h13, 8'h0b, 8'h09, 8'hff, 8'h0d, 8'h07, 8'hf7, 8'hff, 8'h12, 8'hee, 8'h0a, 8'h13, 8'hf0, 8'hfe, 8'h0e, 8'h13, 8'hf9, 8'hff, 8'hec, 8'h01, 8'h10, 8'h0c, 8'h07, 8'hfd, 8'h04, 8'h12, 8'hee, 8'h05, 8'hfb, 8'h11, 8'hfb, 8'h0b, 8'hf6, 8'hfb, 8'h14, 8'h03, 8'h07, 8'hf9};
assign weight_matrix[33] = {8'h13, 8'hfd, 8'h0f, 8'h10, 8'h12, 8'hff, 8'hfd, 8'heb, 8'h02, 8'h0b, 8'hf0, 8'h02, 8'h06, 8'h11, 8'h02, 8'hf6, 8'h06, 8'h12, 8'hec, 8'h11, 8'h00, 8'hfd, 8'h11, 8'hfa, 8'hfc, 8'h0b, 8'hf1, 8'h07, 8'heb, 8'h04, 8'h05, 8'hf1, 8'hf7, 8'hf0, 8'h18, 8'h14, 8'he7, 8'h0b, 8'hf5, 8'hef, 8'h15, 8'hf3, 8'h0c, 8'hfe, 8'h0c, 8'h04, 8'h00, 8'hf4, 8'hfc, 8'h16, 8'h11, 8'hef, 8'hfe, 8'hf9, 8'h02, 8'hfc, 8'hfb, 8'hf9, 8'hf9, 8'h12, 8'h09, 8'h0a, 8'h04, 8'h0e};
assign weight_matrix[34] = {8'h06, 8'hef, 8'h13, 8'h05, 8'hff, 8'h16, 8'h1a, 8'hf4, 8'h07, 8'h06, 8'h05, 8'hf1, 8'h19, 8'h08, 8'hf2, 8'hf7, 8'hf8, 8'hfd, 8'h00, 8'hfc, 8'h0f, 8'h03, 8'heb, 8'h16, 8'he6, 8'hf0, 8'hf5, 8'hf5, 8'hf8, 8'h11, 8'hf1, 8'h14, 8'heb, 8'hfe, 8'h14, 8'hf0, 8'heb, 8'hfd, 8'hff, 8'hf7, 8'h11, 8'h0a, 8'h02, 8'hfa, 8'h09, 8'hff, 8'hf2, 8'h03, 8'hfc, 8'h04, 8'hf2, 8'h02, 8'h10, 8'h12, 8'h0b, 8'h0b, 8'hee, 8'h03, 8'he5, 8'h0b, 8'hfa, 8'h08, 8'he8, 8'h02};
assign weight_matrix[35] = {8'hf9, 8'hde, 8'h0d, 8'hf7, 8'hf6, 8'hef, 8'h0d, 8'hf6, 8'h1c, 8'hf0, 8'he9, 8'h09, 8'h0c, 8'h0d, 8'hf6, 8'hfa, 8'h10, 8'hef, 8'h10, 8'h0d, 8'hf4, 8'hef, 8'hf4, 8'hf9, 8'hfa, 8'he9, 8'h05, 8'h13, 8'h06, 8'h07, 8'hfb, 8'h10, 8'hfc, 8'h13, 8'hf8, 8'hf6, 8'h0d, 8'hf2, 8'hfe, 8'hf4, 8'h06, 8'he7, 8'hee, 8'h04, 8'h14, 8'h02, 8'hea, 8'he6, 8'h0d, 8'hf7, 8'h08, 8'h0e, 8'h02, 8'hea, 8'h01, 8'hf0, 8'h08, 8'hf9, 8'he9, 8'he8, 8'hf9, 8'he2, 8'hf9, 8'h12};
assign weight_matrix[36] = {8'h01, 8'h0f, 8'hfc, 8'hff, 8'hfe, 8'hf5, 8'h15, 8'hf0, 8'h00, 8'hf9, 8'hef, 8'hf4, 8'hf7, 8'h0e, 8'h0c, 8'he7, 8'hed, 8'h01, 8'h0b, 8'hf7, 8'h02, 8'hf8, 8'h00, 8'hfc, 8'h10, 8'hfd, 8'hf7, 8'h00, 8'hf0, 8'hef, 8'h05, 8'h02, 8'hfe, 8'h14, 8'hf1, 8'hec, 8'hee, 8'he9, 8'heb, 8'hf9, 8'h12, 8'h0f, 8'hfc, 8'h0a, 8'hff, 8'hf1, 8'h0e, 8'h05, 8'h0a, 8'hf4, 8'h0b, 8'h13, 8'h0e, 8'hfa, 8'hf0, 8'h0d, 8'h08, 8'h0a, 8'hfb, 8'heb, 8'hf5, 8'h0d, 8'h02, 8'h02};
assign weight_matrix[37] = {8'hfc, 8'hed, 8'hf8, 8'h0b, 8'hf4, 8'h0d, 8'h09, 8'hf7, 8'h0e, 8'hf0, 8'hf7, 8'hf3, 8'hfe, 8'he9, 8'h06, 8'h13, 8'h13, 8'h08, 8'hef, 8'hfa, 8'hf8, 8'h01, 8'h0e, 8'h09, 8'hfa, 8'hfd, 8'h11, 8'hf0, 8'h06, 8'h0f, 8'h01, 8'h13, 8'h07, 8'hf9, 8'h02, 8'h0e, 8'hfd, 8'h12, 8'hf6, 8'h14, 8'h06, 8'hfc, 8'h01, 8'hf9, 8'hf5, 8'h0c, 8'he8, 8'heb, 8'h06, 8'hf7, 8'hff, 8'h17, 8'he9, 8'hed, 8'heb, 8'h11, 8'hfc, 8'h08, 8'hf3, 8'h06, 8'hec, 8'hf4, 8'h09, 8'h17};
assign weight_matrix[38] = {8'h11, 8'h0e, 8'h04, 8'hff, 8'hf0, 8'h12, 8'hfc, 8'hfb, 8'hfd, 8'h02, 8'h0b, 8'h13, 8'hea, 8'h00, 8'h00, 8'hf8, 8'h15, 8'h03, 8'h08, 8'h0a, 8'h11, 8'h14, 8'h0c, 8'h0d, 8'hf3, 8'hfd, 8'h0e, 8'hea, 8'hec, 8'h13, 8'hf9, 8'h07, 8'h07, 8'hef, 8'h0a, 8'h0f, 8'hee, 8'hf0, 8'hfc, 8'hf9, 8'h0f, 8'hf2, 8'h10, 8'h11, 8'hfb, 8'h14, 8'hf0, 8'hee, 8'h06, 8'h03, 8'h01, 8'h08, 8'h0a, 8'h12, 8'hf0, 8'hfe, 8'h01, 8'h15, 8'h0d, 8'h0d, 8'hee, 8'hf4, 8'h14, 8'h05};
assign weight_matrix[39] = {8'hee, 8'h01, 8'h0e, 8'hff, 8'h01, 8'heb, 8'h0b, 8'hf7, 8'hf1, 8'h0e, 8'h0c, 8'hf8, 8'h0b, 8'h01, 8'h10, 8'hf7, 8'hf7, 8'hea, 8'hfa, 8'h0b, 8'h14, 8'h0f, 8'h15, 8'hf6, 8'h04, 8'h15, 8'hf9, 8'h08, 8'h13, 8'h12, 8'hf7, 8'h15, 8'hf6, 8'hea, 8'h10, 8'h01, 8'h0e, 8'h0f, 8'hf2, 8'h00, 8'h0a, 8'h14, 8'h11, 8'h03, 8'h0e, 8'h15, 8'h04, 8'h13, 8'hef, 8'hea, 8'hea, 8'hec, 8'hf1, 8'hea, 8'hec, 8'hfa, 8'hfa, 8'h08, 8'h07, 8'h12, 8'hf1, 8'h0a, 8'h08, 8'hff};
assign weight_matrix[40] = {8'hf1, 8'h0b, 8'h0e, 8'hfe, 8'hf0, 8'hf4, 8'hf5, 8'h03, 8'hf1, 8'h07, 8'h02, 8'hfe, 8'h08, 8'h02, 8'h04, 8'h07, 8'h11, 8'h11, 8'h02, 8'h16, 8'h06, 8'h07, 8'h01, 8'h01, 8'hfa, 8'hef, 8'hfa, 8'hf4, 8'h00, 8'h0a, 8'h13, 8'hf7, 8'h07, 8'hed, 8'h0e, 8'hf2, 8'h0d, 8'h13, 8'hfd, 8'h08, 8'h0a, 8'hed, 8'h0e, 8'hee, 8'heb, 8'h12, 8'h0c, 8'h0c, 8'hf5, 8'hfb, 8'h0e, 8'h0b, 8'hfc, 8'hee, 8'hed, 8'h14, 8'h0c, 8'hfa, 8'hfa, 8'hfd, 8'hec, 8'hee, 8'h0e, 8'hec};
assign weight_matrix[41] = {8'h0a, 8'hf3, 8'h06, 8'h01, 8'hf2, 8'hfc, 8'h0e, 8'h0d, 8'h0c, 8'hf7, 8'h08, 8'hfb, 8'hff, 8'hec, 8'h08, 8'hef, 8'h0d, 8'h02, 8'h0e, 8'h07, 8'h10, 8'h11, 8'h0d, 8'hfb, 8'h01, 8'hea, 8'hed, 8'he8, 8'hea, 8'hfd, 8'hf4, 8'heb, 8'hf1, 8'h0c, 8'h0e, 8'he8, 8'h09, 8'hf2, 8'h11, 8'hf9, 8'h11, 8'hfe, 8'h0a, 8'h07, 8'hee, 8'hf2, 8'h03, 8'h11, 8'h06, 8'h00, 8'hef, 8'he6, 8'h13, 8'h0a, 8'h04, 8'hfc, 8'h12, 8'hf0, 8'hf2, 8'hf1, 8'h04, 8'h0d, 8'h0d, 8'hf1};
assign weight_matrix[42] = {8'he3, 8'h02, 8'h0b, 8'hf9, 8'h04, 8'hfc, 8'hec, 8'he6, 8'hed, 8'h21, 8'h09, 8'h06, 8'hf3, 8'h03, 8'h12, 8'h01, 8'h08, 8'h03, 8'hf0, 8'hfc, 8'h02, 8'hed, 8'h0d, 8'h19, 8'h06, 8'h08, 8'hea, 8'hee, 8'hf7, 8'h13, 8'h07, 8'hd8, 8'hf8, 8'hee, 8'hfb, 8'he8, 8'hf2, 8'hf3, 8'h0e, 8'h19, 8'h00, 8'h03, 8'he7, 8'h00, 8'h17, 8'hf7, 8'hfa, 8'hff, 8'hec, 8'hf2, 8'h18, 8'h00, 8'hf1, 8'h12, 8'h2a, 8'hee, 8'h0e, 8'h23, 8'h09, 8'he7, 8'hf9, 8'h02, 8'hf6, 8'he5};
assign weight_matrix[43] = {8'h06, 8'h04, 8'hfb, 8'h07, 8'h05, 8'hf4, 8'he4, 8'hfc, 8'hff, 8'h0d, 8'h0b, 8'hf5, 8'h00, 8'he9, 8'hf2, 8'hfb, 8'hea, 8'h0c, 8'hf6, 8'heb, 8'hfc, 8'h00, 8'he7, 8'hf6, 8'hf1, 8'h03, 8'hfb, 8'h04, 8'hf5, 8'h03, 8'hf4, 8'h07, 8'h01, 8'hf5, 8'hf1, 8'he9, 8'hf4, 8'he8, 8'hfb, 8'h02, 8'hfd, 8'hf3, 8'hf0, 8'h04, 8'hfa, 8'hf9, 8'hfc, 8'hf9, 8'hf2, 8'hf4, 8'hf7, 8'hfc, 8'hf3, 8'hfe, 8'h02, 8'he8, 8'hf8, 8'h0e, 8'hee, 8'hfa, 8'h07, 8'h0b, 8'h09, 8'h0a};
assign weight_matrix[44] = {8'h12, 8'h03, 8'hfe, 8'hfb, 8'h0f, 8'h05, 8'hf6, 8'h10, 8'hfe, 8'h07, 8'h06, 8'hf6, 8'h07, 8'hf5, 8'h16, 8'h0d, 8'hf1, 8'h04, 8'hed, 8'hef, 8'h07, 8'h0a, 8'hf0, 8'h0b, 8'h00, 8'h0a, 8'hf5, 8'hf7, 8'h09, 8'h0b, 8'hf4, 8'h08, 8'h10, 8'hf6, 8'h0a, 8'h11, 8'h06, 8'h07, 8'hfc, 8'h13, 8'hfc, 8'hea, 8'hf0, 8'h15, 8'hfa, 8'h12, 8'h09, 8'hfd, 8'h14, 8'hf0, 8'h11, 8'hea, 8'hea, 8'h01, 8'hfd, 8'h0c, 8'hfc, 8'hfb, 8'hf5, 8'h04, 8'h15, 8'h0e, 8'hf8, 8'h0e};
assign weight_matrix[45] = {8'h17, 8'hfc, 8'h05, 8'hec, 8'he7, 8'hef, 8'hee, 8'h06, 8'h07, 8'h17, 8'hf3, 8'h16, 8'hed, 8'he9, 8'hf3, 8'hfe, 8'h0f, 8'h11, 8'h05, 8'he9, 8'h0a, 8'hf9, 8'hec, 8'h09, 8'hf0, 8'hd5, 8'h0f, 8'h07, 8'h01, 8'hf8, 8'h07, 8'he9, 8'hed, 8'h01, 8'h11, 8'hee, 8'h0b, 8'hf9, 8'hff, 8'h01, 8'hfc, 8'h0d, 8'hf0, 8'hf0, 8'h01, 8'hf5, 8'hfd, 8'h09, 8'hef, 8'hfe, 8'hf8, 8'hf7, 8'h08, 8'h0e, 8'h05, 8'h00, 8'h11, 8'hfe, 8'hd3, 8'h0d, 8'hed, 8'h10, 8'h11, 8'hfb};
assign weight_matrix[46] = {8'h0d, 8'hf2, 8'hef, 8'h16, 8'h11, 8'h13, 8'hfb, 8'hfe, 8'h07, 8'h06, 8'hf5, 8'hfd, 8'hf8, 8'h03, 8'h07, 8'hf3, 8'h02, 8'h13, 8'h07, 8'h0b, 8'h02, 8'h10, 8'hee, 8'h06, 8'hee, 8'h02, 8'h07, 8'h14, 8'h11, 8'h02, 8'hf9, 8'h13, 8'hf3, 8'hf5, 8'hed, 8'hfd, 8'hf7, 8'h04, 8'h05, 8'hea, 8'hfd, 8'h14, 8'hf9, 8'hec, 8'hf7, 8'h16, 8'hea, 8'h02, 8'h0a, 8'h02, 8'hf8, 8'hfe, 8'hf2, 8'h08, 8'hf3, 8'h0a, 8'hea, 8'h13, 8'h16, 8'h0a, 8'hf7, 8'hfb, 8'hfc, 8'hf2};
assign weight_matrix[47] = {8'hf4, 8'hf2, 8'hea, 8'hf2, 8'h09, 8'hf3, 8'heb, 8'hff, 8'hfe, 8'hf3, 8'h0b, 8'h09, 8'h16, 8'hf9, 8'h08, 8'h03, 8'h09, 8'hf4, 8'h0a, 8'hf3, 8'h0e, 8'hf6, 8'hf7, 8'h0f, 8'h0a, 8'hf2, 8'h16, 8'hfa, 8'h16, 8'h00, 8'hf6, 8'h09, 8'h08, 8'hf5, 8'h16, 8'h00, 8'hea, 8'h0f, 8'hf6, 8'h15, 8'h08, 8'h05, 8'hfb, 8'hfc, 8'h0d, 8'h12, 8'h10, 8'h03, 8'hf2, 8'h0c, 8'h02, 8'h03, 8'h16, 8'hec, 8'h11, 8'h09, 8'h00, 8'h00, 8'h0c, 8'hed, 8'h0c, 8'h04, 8'h02, 8'h13};
assign weight_matrix[48] = {8'hf5, 8'h0a, 8'h0a, 8'h0f, 8'h02, 8'heb, 8'h0d, 8'hee, 8'he7, 8'h03, 8'h12, 8'hf6, 8'he8, 8'hf4, 8'h0c, 8'hf8, 8'hed, 8'he7, 8'hf0, 8'hfd, 8'h0a, 8'hf8, 8'hec, 8'h09, 8'hf1, 8'hfb, 8'heb, 8'hf7, 8'hf5, 8'hfc, 8'he4, 8'h10, 8'h0e, 8'hf0, 8'h10, 8'hed, 8'h0c, 8'h0a, 8'h0a, 8'he5, 8'h11, 8'hf4, 8'hfd, 8'h14, 8'hf6, 8'h01, 8'hf3, 8'hf4, 8'h08, 8'hf0, 8'h06, 8'h0f, 8'hf5, 8'h12, 8'h0a, 8'hee, 8'hed, 8'h09, 8'h1a, 8'he6, 8'hee, 8'hf5, 8'hfd, 8'h06};
assign weight_matrix[49] = {8'hef, 8'hfe, 8'h0e, 8'h00, 8'hf7, 8'h03, 8'h00, 8'hf9, 8'hec, 8'h08, 8'h14, 8'h03, 8'h16, 8'hfa, 8'h0d, 8'h16, 8'hed, 8'h12, 8'h01, 8'h15, 8'h01, 8'hf4, 8'h05, 8'h04, 8'hf6, 8'h13, 8'h10, 8'h0e, 8'h00, 8'hfa, 8'hfe, 8'h02, 8'h01, 8'hf0, 8'h01, 8'hff, 8'h0f, 8'hf1, 8'hf2, 8'hec, 8'h0a, 8'hfb, 8'heb, 8'hfd, 8'h12, 8'hf7, 8'hec, 8'hff, 8'hf5, 8'hf2, 8'h12, 8'hf1, 8'h00, 8'hfa, 8'hf5, 8'hf4, 8'h0d, 8'h00, 8'hfa, 8'hf4, 8'h03, 8'hfe, 8'h0d, 8'h0a};
assign weight_matrix[50] = {8'h0e, 8'he9, 8'heb, 8'h09, 8'he9, 8'hfb, 8'hf1, 8'h06, 8'hfa, 8'hf3, 8'hf6, 8'heb, 8'h02, 8'h05, 8'h06, 8'heb, 8'h08, 8'h01, 8'hff, 8'h09, 8'hfe, 8'hec, 8'h12, 8'h10, 8'h07, 8'he4, 8'h03, 8'h0f, 8'hfb, 8'heb, 8'hee, 8'h10, 8'he6, 8'hfd, 8'h0a, 8'hf7, 8'h04, 8'hf6, 8'heb, 8'hea, 8'hf4, 8'hf0, 8'hf0, 8'h0b, 8'h09, 8'h0b, 8'h05, 8'hec, 8'hfa, 8'h00, 8'h03, 8'hed, 8'hf7, 8'h07, 8'h08, 8'h01, 8'hff, 8'h0c, 8'h03, 8'hea, 8'hf9, 8'h05, 8'h0b, 8'h0c};
assign weight_matrix[51] = {8'h05, 8'h0d, 8'heb, 8'h19, 8'he9, 8'h18, 8'h0b, 8'h04, 8'h08, 8'hdd, 8'h1a, 8'hf3, 8'h0d, 8'hfd, 8'h08, 8'h04, 8'hf1, 8'hef, 8'he5, 8'hee, 8'h0c, 8'hfa, 8'h07, 8'hf3, 8'hf4, 8'h06, 8'hf9, 8'hf8, 8'hf4, 8'hf1, 8'hfc, 8'heb, 8'hdb, 8'h08, 8'hfb, 8'h0c, 8'hf2, 8'h00, 8'hf0, 8'h13, 8'h11, 8'h00, 8'hff, 8'h0e, 8'h07, 8'hf0, 8'h0f, 8'hf9, 8'hf9, 8'hf9, 8'hf5, 8'hfc, 8'h18, 8'h12, 8'hf7, 8'hf5, 8'hec, 8'h1e, 8'h00, 8'hf6, 8'hfc, 8'hf1, 8'hed, 8'hf0};
assign weight_matrix[52] = {8'hf8, 8'hf2, 8'hfd, 8'h0d, 8'hf0, 8'hf5, 8'hf3, 8'hfd, 8'hf3, 8'hf6, 8'hf3, 8'h09, 8'hed, 8'h08, 8'h08, 8'h0e, 8'h0c, 8'hed, 8'hf6, 8'hf7, 8'hf9, 8'hec, 8'hfc, 8'hf5, 8'h02, 8'hf9, 8'h0a, 8'h09, 8'hf5, 8'hef, 8'hee, 8'h11, 8'hfc, 8'hfd, 8'heb, 8'h01, 8'hf0, 8'h07, 8'hfc, 8'h0e, 8'h0d, 8'h08, 8'h0a, 8'h0d, 8'hfc, 8'hfa, 8'hff, 8'h0c, 8'hf5, 8'hf4, 8'h0a, 8'hfe, 8'hea, 8'hfb, 8'h02, 8'hee, 8'heb, 8'h00, 8'h15, 8'h07, 8'hfa, 8'h0c, 8'hff, 8'hfa};
assign weight_matrix[53] = {8'h11, 8'h05, 8'hfc, 8'hfd, 8'h08, 8'h04, 8'h0a, 8'h0e, 8'h0c, 8'hf1, 8'hfb, 8'hed, 8'hff, 8'h10, 8'heb, 8'h13, 8'h01, 8'hfc, 8'h0f, 8'h0d, 8'h0b, 8'he9, 8'hfa, 8'hf3, 8'h07, 8'hfa, 8'hf3, 8'h11, 8'hfc, 8'hed, 8'he9, 8'h08, 8'hf1, 8'h03, 8'hf0, 8'hf1, 8'h06, 8'h02, 8'h01, 8'hf2, 8'hf8, 8'hf8, 8'hed, 8'hfe, 8'h07, 8'he9, 8'hf0, 8'hf4, 8'hef, 8'h00, 8'hfa, 8'hf0, 8'hf8, 8'hf5, 8'hf4, 8'hf2, 8'h04, 8'hf6, 8'heb, 8'hf8, 8'h0f, 8'hfb, 8'hfe, 8'h12};
assign weight_matrix[54] = {8'h03, 8'h07, 8'hf9, 8'h0a, 8'h0e, 8'h11, 8'hf8, 8'h13, 8'h06, 8'h0b, 8'hff, 8'hff, 8'h00, 8'hff, 8'hf2, 8'hef, 8'h06, 8'h03, 8'h0a, 8'hec, 8'hf2, 8'h02, 8'h08, 8'hfa, 8'heb, 8'hfc, 8'h08, 8'hfe, 8'h0d, 8'hff, 8'hfd, 8'h06, 8'hff, 8'he9, 8'hf5, 8'hf9, 8'h01, 8'hea, 8'hfe, 8'h0a, 8'h05, 8'hf2, 8'hf2, 8'h02, 8'h08, 8'hec, 8'h09, 8'h0c, 8'hec, 8'hfc, 8'h0a, 8'hfe, 8'he9, 8'hef, 8'h12, 8'hf0, 8'hf1, 8'h06, 8'hf7, 8'hf2, 8'h0a, 8'hf9, 8'h08, 8'hf7};
assign weight_matrix[55] = {8'hfd, 8'h04, 8'h03, 8'hfb, 8'h01, 8'h17, 8'h09, 8'heb, 8'h0c, 8'h00, 8'hfa, 8'h11, 8'h15, 8'h10, 8'hfb, 8'hec, 8'h14, 8'h0c, 8'h14, 8'h08, 8'h0f, 8'hf3, 8'h01, 8'h06, 8'h12, 8'hef, 8'h13, 8'he9, 8'hf9, 8'h11, 8'hf5, 8'h15, 8'h11, 8'h03, 8'h08, 8'hee, 8'hf5, 8'h05, 8'h10, 8'hf0, 8'hed, 8'h0a, 8'h0c, 8'hde, 8'hf3, 8'hee, 8'hfa, 8'hf7, 8'h00, 8'hf8, 8'hf7, 8'hf8, 8'hfc, 8'h08, 8'h13, 8'hfc, 8'heb, 8'hee, 8'hfa, 8'h00, 8'hf9, 8'hec, 8'h01, 8'hf5};
assign weight_matrix[56] = {8'h06, 8'h0b, 8'h10, 8'hf8, 8'h01, 8'h08, 8'h0d, 8'h0a, 8'h00, 8'hff, 8'h02, 8'hfc, 8'h00, 8'hf8, 8'hf4, 8'h07, 8'hf6, 8'h05, 8'hfb, 8'hef, 8'hff, 8'hfa, 8'h0b, 8'h04, 8'hfb, 8'h10, 8'hf6, 8'hff, 8'hec, 8'h13, 8'hfb, 8'h0d, 8'hec, 8'hf9, 8'hf6, 8'h0b, 8'hf6, 8'hf9, 8'h14, 8'h10, 8'h0b, 8'hf7, 8'hfb, 8'h16, 8'h0b, 8'hfb, 8'hf7, 8'h06, 8'hfe, 8'h0b, 8'hf7, 8'h18, 8'hf7, 8'h00, 8'hf3, 8'h07, 8'h07, 8'h18, 8'he2, 8'hee, 8'hff, 8'hfa, 8'hed, 8'hf0};
assign weight_matrix[57] = {8'hf8, 8'h2b, 8'h0c, 8'h0b, 8'h02, 8'he9, 8'he4, 8'h12, 8'hf3, 8'h18, 8'h07, 8'hf8, 8'hfa, 8'h05, 8'hf8, 8'he9, 8'hfe, 8'hfa, 8'he7, 8'hec, 8'hf6, 8'he7, 8'hf4, 8'hfc, 8'h03, 8'hee, 8'hea, 8'hed, 8'h09, 8'h29, 8'hef, 8'heb, 8'hfe, 8'hf0, 8'hfb, 8'h17, 8'hed, 8'hfe, 8'h19, 8'h18, 8'h23, 8'h18, 8'h0a, 8'h05, 8'hed, 8'h0d, 8'h03, 8'h25, 8'hf0, 8'h1b, 8'h00, 8'hfc, 8'hfd, 8'hec, 8'hee, 8'h03, 8'h14, 8'h24, 8'h14, 8'hf7, 8'hf7, 8'h04, 8'he4, 8'hdc};
assign weight_matrix[58] = {8'hd0, 8'h02, 8'h10, 8'h06, 8'h21, 8'h1a, 8'h05, 8'hff, 8'hde, 8'h22, 8'h0c, 8'hee, 8'hf8, 8'hed, 8'heb, 8'h06, 8'h08, 8'hf3, 8'he6, 8'h04, 8'hff, 8'he4, 8'hef, 8'h41, 8'hfd, 8'h05, 8'h09, 8'hec, 8'h0a, 8'h2c, 8'hf2, 8'hbb, 8'h25, 8'heb, 8'he5, 8'hf1, 8'h06, 8'hf5, 8'h09, 8'h13, 8'h0b, 8'h16, 8'h18, 8'hec, 8'h25, 8'h20, 8'he8, 8'hee, 8'h06, 8'h0d, 8'h20, 8'hef, 8'hf3, 8'h07, 8'h30, 8'h0b, 8'he8, 8'h55, 8'h0a, 8'h0c, 8'hf0, 8'h44, 8'hc7, 8'hc9};
assign weight_matrix[59] = {8'h07, 8'hf7, 8'h08, 8'h13, 8'hed, 8'h0b, 8'h0d, 8'hf0, 8'heb, 8'h01, 8'he9, 8'hf6, 8'h14, 8'hf8, 8'h01, 8'h04, 8'h04, 8'h09, 8'h06, 8'h0d, 8'h0a, 8'h05, 8'hf6, 8'hfd, 8'h07, 8'he6, 8'h01, 8'h12, 8'hf0, 8'hff, 8'hec, 8'h0a, 8'hfe, 8'hf0, 8'hf7, 8'hed, 8'h0d, 8'h06, 8'h03, 8'hef, 8'h0f, 8'hfe, 8'h06, 8'hed, 8'h0b, 8'hed, 8'h05, 8'hf8, 8'hed, 8'hff, 8'hec, 8'h0a, 8'hfd, 8'h09, 8'h06, 8'h08, 8'h0d, 8'hec, 8'h04, 8'h11, 8'h0c, 8'hfd, 8'h1d, 8'h15};
assign weight_matrix[60] = {8'hff, 8'hf0, 8'h0c, 8'h13, 8'hfe, 8'hf4, 8'hf2, 8'hfd, 8'h08, 8'h0a, 8'hf5, 8'hf0, 8'hfa, 8'h0b, 8'h16, 8'h0d, 8'hfa, 8'hf8, 8'h0e, 8'h16, 8'hfb, 8'hf0, 8'h04, 8'h16, 8'hef, 8'hff, 8'h05, 8'h05, 8'hf7, 8'h08, 8'hfd, 8'hf6, 8'h07, 8'h0f, 8'h0e, 8'h06, 8'hf8, 8'h02, 8'h03, 8'h14, 8'hf3, 8'hf9, 8'h0d, 8'h05, 8'hf4, 8'hf8, 8'hf2, 8'h0a, 8'h10, 8'h13, 8'h04, 8'hf7, 8'hfd, 8'h0b, 8'h10, 8'hf4, 8'h06, 8'h03, 8'hea, 8'hf2, 8'h0a, 8'hfc, 8'h12, 8'hfd};
assign weight_matrix[61] = {8'hfa, 8'h14, 8'hff, 8'hf7, 8'h0a, 8'h00, 8'hf5, 8'hf3, 8'h05, 8'hef, 8'hf0, 8'hfd, 8'h02, 8'h0b, 8'hfb, 8'h02, 8'he7, 8'he8, 8'h02, 8'h04, 8'heb, 8'h06, 8'h03, 8'hfc, 8'hf4, 8'hf7, 8'h03, 8'hf2, 8'h08, 8'h05, 8'hec, 8'hfb, 8'hf2, 8'hfc, 8'hf7, 8'hf3, 8'hf6, 8'h11, 8'hec, 8'h02, 8'hee, 8'h0a, 8'hfe, 8'hfa, 8'hed, 8'hf3, 8'hf3, 8'h03, 8'hf0, 8'hf9, 8'h09, 8'heb, 8'h08, 8'hfa, 8'hf6, 8'h0b, 8'h0b, 8'h03, 8'hf0, 8'hec, 8'hfb, 8'h15, 8'h03, 8'h12};
assign weight_matrix[62] = {8'hf1, 8'h04, 8'hf8, 8'h0c, 8'hed, 8'hed, 8'h15, 8'hff, 8'hfc, 8'hf7, 8'h0e, 8'h08, 8'hf5, 8'h13, 8'h0a, 8'hf9, 8'h13, 8'hf0, 8'h02, 8'hee, 8'h0b, 8'h02, 8'h01, 8'h02, 8'h0c, 8'h14, 8'h0d, 8'h0a, 8'h02, 8'hf3, 8'h05, 8'h01, 8'h06, 8'h10, 8'hfc, 8'h02, 8'hfe, 8'hec, 8'hf1, 8'h0a, 8'hfa, 8'hed, 8'hf1, 8'hf4, 8'h09, 8'hfe, 8'hf5, 8'hf6, 8'hf8, 8'hfb, 8'h02, 8'hee, 8'h0d, 8'h15, 8'h16, 8'h16, 8'hfb, 8'h02, 8'h08, 8'hf9, 8'h12, 8'h03, 8'hf1, 8'hf1};
assign weight_matrix[63] = {8'hff, 8'h0e, 8'h12, 8'hed, 8'hfc, 8'hf3, 8'heb, 8'h0e, 8'hee, 8'hee, 8'hef, 8'hf0, 8'h16, 8'h07, 8'h15, 8'hfa, 8'h0a, 8'hfa, 8'hed, 8'hf6, 8'hf2, 8'h03, 8'h06, 8'hf3, 8'hf8, 8'h08, 8'h10, 8'h16, 8'hef, 8'h0e, 8'h03, 8'h03, 8'hfd, 8'h01, 8'h12, 8'hf5, 8'h05, 8'h02, 8'hf4, 8'h16, 8'hf5, 8'hf9, 8'h00, 8'hf0, 8'hf6, 8'hfa, 8'h0d, 8'hed, 8'heb, 8'h13, 8'h0e, 8'hfc, 8'h0a, 8'h03, 8'h0e, 8'h01, 8'hea, 8'hf8, 8'hfd, 8'hec, 8'hff, 8'hee, 8'hfc, 8'h00};
assign weight_matrix[64] = {8'h05, 8'hea, 8'hf3, 8'hf0, 8'h04, 8'h01, 8'hf6, 8'hf3, 8'hfa, 8'h09, 8'h0b, 8'h06, 8'h00, 8'h07, 8'hf8, 8'hf2, 8'hf2, 8'h07, 8'h0b, 8'hec, 8'hfe, 8'hea, 8'h07, 8'hf5, 8'hed, 8'h0c, 8'he9, 8'hea, 8'h14, 8'h07, 8'hfd, 8'hf0, 8'h05, 8'hf9, 8'h0f, 8'hfd, 8'h06, 8'hfd, 8'hf6, 8'hff, 8'he9, 8'hf0, 8'h0e, 8'h0c, 8'h0a, 8'hf1, 8'hee, 8'hff, 8'hfb, 8'h0a, 8'hf6, 8'hfe, 8'hfe, 8'h10, 8'hef, 8'h01, 8'hff, 8'hfe, 8'hdd, 8'h0a, 8'hfe, 8'hf9, 8'hfa, 8'h0b};
assign weight_matrix[65] = {8'he4, 8'h0c, 8'hfb, 8'h0f, 8'h15, 8'hea, 8'hf4, 8'h0f, 8'h0a, 8'hfd, 8'h03, 8'hff, 8'he8, 8'he9, 8'hfd, 8'hed, 8'h15, 8'h07, 8'hef, 8'h04, 8'h07, 8'h08, 8'h07, 8'h11, 8'hec, 8'h08, 8'h14, 8'hf8, 8'h15, 8'h07, 8'hf9, 8'heb, 8'hf3, 8'hf4, 8'h0f, 8'hea, 8'h11, 8'h09, 8'h11, 8'h00, 8'h0e, 8'h17, 8'h11, 8'h12, 8'h07, 8'h11, 8'h07, 8'hee, 8'h05, 8'hf8, 8'h04, 8'h0f, 8'hf1, 8'hf5, 8'h03, 8'hef, 8'h12, 8'h0e, 8'h19, 8'h0b, 8'hf1, 8'h15, 8'hf1, 8'h08};
assign weight_matrix[66] = {8'h0d, 8'hff, 8'hf5, 8'h0c, 8'h0a, 8'h01, 8'hf8, 8'hec, 8'h07, 8'hf4, 8'h0e, 8'hf4, 8'h12, 8'hf7, 8'h00, 8'h08, 8'h02, 8'hf4, 8'hfb, 8'hfc, 8'hf3, 8'hf4, 8'h0f, 8'h0f, 8'hf7, 8'hef, 8'h0a, 8'hfb, 8'hf5, 8'hee, 8'heb, 8'hfb, 8'he8, 8'hf8, 8'hee, 8'h0b, 8'h15, 8'hfc, 8'hf7, 8'hfb, 8'hf2, 8'hfd, 8'h0d, 8'hf9, 8'h0e, 8'h0c, 8'hf1, 8'h04, 8'heb, 8'hf7, 8'hef, 8'hfa, 8'h01, 8'h0b, 8'hff, 8'h02, 8'hf0, 8'hf1, 8'he7, 8'h10, 8'h04, 8'hf7, 8'h03, 8'hf1};
assign weight_matrix[67] = {8'hfa, 8'hf6, 8'h09, 8'hf7, 8'h0d, 8'h11, 8'hec, 8'hef, 8'hfa, 8'h1c, 8'h07, 8'hfd, 8'h06, 8'hf5, 8'h02, 8'hfa, 8'hff, 8'h0e, 8'h15, 8'h09, 8'hf1, 8'hef, 8'hf1, 8'he7, 8'h0e, 8'hec, 8'hf7, 8'hf0, 8'hf3, 8'hfa, 8'hfb, 8'h0a, 8'he9, 8'hff, 8'h15, 8'h0d, 8'h0b, 8'hfa, 8'h02, 8'hfe, 8'h01, 8'h03, 8'hff, 8'hef, 8'hf1, 8'h10, 8'hf2, 8'h0a, 8'h0a, 8'hf1, 8'h08, 8'h08, 8'h0b, 8'he8, 8'hfa, 8'h11, 8'h00, 8'hf2, 8'h06, 8'h0f, 8'hfc, 8'hec, 8'h12, 8'h17};
assign weight_matrix[68] = {8'he2, 8'hf1, 8'h15, 8'h07, 8'h14, 8'h03, 8'h12, 8'hec, 8'he3, 8'h30, 8'he5, 8'h18, 8'hec, 8'h0d, 8'h05, 8'h07, 8'h1c, 8'h11, 8'h0c, 8'he2, 8'h06, 8'h01, 8'h1a, 8'h30, 8'hf4, 8'hda, 8'h04, 8'hf1, 8'hf4, 8'h36, 8'hfc, 8'hde, 8'h4f, 8'hfc, 8'h0c, 8'he6, 8'h07, 8'hf6, 8'h0b, 8'h0b, 8'h18, 8'h1d, 8'hfd, 8'hcf, 8'hfe, 8'h15, 8'hef, 8'hf9, 8'h06, 8'h08, 8'h1f, 8'hf8, 8'hf0, 8'hec, 8'h20, 8'h05, 8'h03, 8'h18, 8'h12, 8'h07, 8'h09, 8'h1b, 8'he6, 8'h03};
assign weight_matrix[69] = {8'hfd, 8'hf3, 8'hff, 8'h13, 8'h0f, 8'hec, 8'hea, 8'h11, 8'hea, 8'hf3, 8'hf3, 8'hf7, 8'hf9, 8'hec, 8'hfd, 8'hf4, 8'h14, 8'hed, 8'h11, 8'h01, 8'h0d, 8'hed, 8'hea, 8'hf6, 8'hec, 8'h0d, 8'hf5, 8'h0c, 8'h03, 8'heb, 8'hf4, 8'h0e, 8'h0b, 8'h0e, 8'hf1, 8'h14, 8'h00, 8'hec, 8'hf9, 8'h06, 8'hef, 8'hf4, 8'hfb, 8'h0b, 8'hfc, 8'hf2, 8'hfe, 8'h10, 8'h0a, 8'h07, 8'h03, 8'hf9, 8'h09, 8'h00, 8'hf7, 8'hf4, 8'h06, 8'h10, 8'h03, 8'h0a, 8'h0d, 8'hed, 8'h0d, 8'hf4};
assign weight_matrix[70] = {8'hf6, 8'hee, 8'h0f, 8'h0d, 8'hff, 8'hf0, 8'h00, 8'hf2, 8'h0a, 8'hed, 8'h11, 8'he9, 8'h00, 8'h01, 8'hf1, 8'h13, 8'hf3, 8'h00, 8'h0a, 8'h12, 8'hfe, 8'h06, 8'hf4, 8'hfe, 8'hea, 8'hea, 8'hed, 8'hea, 8'hf6, 8'hfe, 8'h01, 8'h16, 8'hee, 8'hff, 8'h03, 8'hfe, 8'hed, 8'hef, 8'hf0, 8'hfe, 8'hf1, 8'hfb, 8'h00, 8'h08, 8'hf8, 8'hea, 8'h0d, 8'hf9, 8'hf6, 8'h0b, 8'hec, 8'hff, 8'h05, 8'h05, 8'h00, 8'hed, 8'h00, 8'hf2, 8'hf5, 8'h08, 8'hf4, 8'hee, 8'h12, 8'h1b};
assign weight_matrix[71] = {8'h07, 8'hf7, 8'hf7, 8'hfb, 8'h04, 8'heb, 8'h04, 8'h01, 8'h04, 8'h1b, 8'h07, 8'h14, 8'h05, 8'hfb, 8'hf4, 8'hfb, 8'h0f, 8'h0f, 8'h02, 8'hf2, 8'hf4, 8'hec, 8'h07, 8'h0e, 8'h09, 8'hf7, 8'hf5, 8'h12, 8'hf8, 8'h14, 8'hf3, 8'h06, 8'h00, 8'hfe, 8'h04, 8'h04, 8'he8, 8'he7, 8'h12, 8'hed, 8'h0d, 8'h18, 8'hf5, 8'hf7, 8'h1a, 8'h1f, 8'h0a, 8'hf3, 8'h08, 8'hef, 8'h01, 8'hfd, 8'hf8, 8'h10, 8'h28, 8'hea, 8'h08, 8'h06, 8'h08, 8'hfe, 8'hef, 8'h05, 8'hef, 8'hec};
assign weight_matrix[72] = {8'h16, 8'hf5, 8'h0d, 8'h01, 8'hf8, 8'h14, 8'h15, 8'h09, 8'h04, 8'heb, 8'h10, 8'h12, 8'h00, 8'hf4, 8'hed, 8'hf4, 8'h0a, 8'hfe, 8'hfa, 8'hfe, 8'h00, 8'h05, 8'hfa, 8'h06, 8'hf3, 8'hf5, 8'hed, 8'hed, 8'h03, 8'h0d, 8'hf1, 8'hfc, 8'hed, 8'hf8, 8'hee, 8'h0b, 8'h0d, 8'h13, 8'h02, 8'h0b, 8'h06, 8'hf0, 8'h05, 8'hf0, 8'h06, 8'h00, 8'hea, 8'h0b, 8'h12, 8'hf2, 8'h11, 8'h0b, 8'h03, 8'hf7, 8'h0e, 8'h08, 8'hff, 8'h03, 8'h08, 8'hf9, 8'h08, 8'h02, 8'h06, 8'hff};
assign weight_matrix[73] = {8'h04, 8'h01, 8'h02, 8'hf1, 8'hf2, 8'hf7, 8'hf6, 8'h0a, 8'h08, 8'h0f, 8'hed, 8'h0d, 8'hea, 8'h05, 8'hf0, 8'h02, 8'hf4, 8'h03, 8'h11, 8'h14, 8'hfa, 8'hf7, 8'hfa, 8'h0d, 8'hec, 8'hf7, 8'hf6, 8'h01, 8'hfa, 8'h05, 8'h11, 8'h06, 8'h09, 8'h0a, 8'hfb, 8'hf4, 8'h14, 8'hf2, 8'h09, 8'h03, 8'h02, 8'h0e, 8'hec, 8'hed, 8'hef, 8'hfe, 8'hf6, 8'hef, 8'hf2, 8'hf1, 8'h05, 8'hfa, 8'hfb, 8'h03, 8'h12, 8'hf8, 8'h15, 8'hf9, 8'heb, 8'hfa, 8'hf1, 8'h0b, 8'h04, 8'hff};
assign weight_matrix[74] = {8'h12, 8'hee, 8'hfa, 8'h0c, 8'hef, 8'heb, 8'h0d, 8'h0f, 8'hfa, 8'hed, 8'h0e, 8'hf3, 8'hec, 8'hf2, 8'hee, 8'h02, 8'h0d, 8'hff, 8'hec, 8'h11, 8'heb, 8'hf9, 8'h0e, 8'hfb, 8'h15, 8'h08, 8'h03, 8'h09, 8'h01, 8'h0e, 8'hf3, 8'h15, 8'hfa, 8'hec, 8'h12, 8'hf4, 8'hef, 8'h03, 8'h12, 8'hf6, 8'h0e, 8'hf9, 8'hf0, 8'h03, 8'h07, 8'h03, 8'h09, 8'hf4, 8'h0b, 8'hf1, 8'h11, 8'h09, 8'h0b, 8'h0d, 8'hf1, 8'hf9, 8'h14, 8'h0c, 8'h0c, 8'hf1, 8'h13, 8'h0d, 8'hf2, 8'hf8};
assign weight_matrix[75] = {8'hea, 8'he0, 8'hec, 8'he6, 8'h12, 8'hed, 8'h0d, 8'hf9, 8'hf8, 8'h22, 8'h07, 8'hef, 8'h0c, 8'h00, 8'hfa, 8'hfa, 8'h08, 8'h0b, 8'hfa, 8'h16, 8'he9, 8'h0e, 8'hf6, 8'hf3, 8'hfa, 8'hfa, 8'hf4, 8'hf2, 8'hed, 8'h0d, 8'hf7, 8'hfe, 8'h17, 8'hf5, 8'hf3, 8'h0e, 8'h03, 8'h14, 8'h06, 8'h18, 8'h0d, 8'h0b, 8'h0e, 8'hf3, 8'hf1, 8'hf7, 8'h06, 8'h04, 8'h16, 8'h12, 8'hed, 8'hf5, 8'h05, 8'h02, 8'h07, 8'hf0, 8'h08, 8'h0a, 8'h13, 8'he7, 8'hf9, 8'h0c, 8'he8, 8'hf2};
assign weight_matrix[76] = {8'hee, 8'h12, 8'h04, 8'hf2, 8'hff, 8'h0b, 8'hff, 8'h12, 8'h0f, 8'hff, 8'h13, 8'h13, 8'hf5, 8'hef, 8'hfb, 8'hf7, 8'hfa, 8'hf1, 8'hea, 8'hea, 8'h15, 8'h00, 8'h09, 8'hf3, 8'h0c, 8'hf5, 8'hf4, 8'hf0, 8'h11, 8'hfa, 8'h02, 8'h07, 8'h0c, 8'h06, 8'hfc, 8'hfb, 8'hfb, 8'h0b, 8'h06, 8'hee, 8'hf6, 8'heb, 8'h15, 8'h04, 8'hff, 8'hfb, 8'hf0, 8'h0c, 8'h16, 8'h0b, 8'h06, 8'h15, 8'hed, 8'h09, 8'hf5, 8'h0f, 8'h05, 8'h04, 8'hf4, 8'h0d, 8'hfc, 8'h14, 8'hea, 8'hfd};
assign weight_matrix[77] = {8'heb, 8'h14, 8'h04, 8'hf8, 8'hf4, 8'hed, 8'h06, 8'h09, 8'h15, 8'hea, 8'h14, 8'hf2, 8'h0f, 8'hf9, 8'heb, 8'h10, 8'he5, 8'h0d, 8'hf2, 8'hf7, 8'h06, 8'h11, 8'hf2, 8'he1, 8'hff, 8'h22, 8'h05, 8'h07, 8'hf2, 8'hee, 8'hef, 8'hfd, 8'he9, 8'he8, 8'h0d, 8'h0f, 8'hfd, 8'hed, 8'hf3, 8'h0c, 8'h08, 8'he5, 8'h0e, 8'h33, 8'h08, 8'he1, 8'h0b, 8'h08, 8'heb, 8'hfb, 8'he3, 8'hf7, 8'hef, 8'hff, 8'he8, 8'h0f, 8'hf8, 8'h20, 8'h02, 8'he7, 8'h02, 8'h06, 8'h00, 8'h13};
assign weight_matrix[78] = {8'h12, 8'hdd, 8'hf6, 8'h03, 8'h0a, 8'hff, 8'he1, 8'h08, 8'h0a, 8'h28, 8'he4, 8'hec, 8'h12, 8'hed, 8'hea, 8'h0a, 8'h0c, 8'h0e, 8'he8, 8'h07, 8'h01, 8'h11, 8'hf5, 8'h05, 8'hfa, 8'hda, 8'h0d, 8'h10, 8'he4, 8'h1a, 8'hea, 8'he5, 8'h2a, 8'hfb, 8'hf8, 8'h10, 8'hf3, 8'hfe, 8'he2, 8'hf7, 8'hff, 8'h10, 8'hf0, 8'hdc, 8'h03, 8'heb, 8'hf5, 8'h0e, 8'hef, 8'h12, 8'h02, 8'hdb, 8'hfa, 8'hed, 8'hfd, 8'hf8, 8'hed, 8'h06, 8'h0c, 8'hf0, 8'hfd, 8'h12, 8'hfd, 8'hfa};
assign weight_matrix[79] = {8'h12, 8'hef, 8'h04, 8'h00, 8'hf1, 8'h0c, 8'h14, 8'h03, 8'hfe, 8'hfc, 8'hfb, 8'hff, 8'hf4, 8'hf9, 8'h16, 8'h11, 8'hfd, 8'h07, 8'hee, 8'h11, 8'h0a, 8'hf9, 8'h04, 8'h0c, 8'hf0, 8'h07, 8'h14, 8'hf2, 8'h16, 8'hfe, 8'h05, 8'hf3, 8'hff, 8'h05, 8'h12, 8'hef, 8'h0b, 8'h06, 8'hfb, 8'h0a, 8'h15, 8'h11, 8'hf3, 8'hf8, 8'h06, 8'h08, 8'h16, 8'h01, 8'h0e, 8'hfc, 8'hf1, 8'h00, 8'hff, 8'hf2, 8'hf4, 8'hf4, 8'h0a, 8'hf1, 8'h0a, 8'hfe, 8'hff, 8'h05, 8'h10, 8'hfe};
assign weight_matrix[80] = {8'hfa, 8'h16, 8'h0c, 8'h04, 8'h18, 8'hea, 8'h01, 8'he8, 8'h0a, 8'hd8, 8'h17, 8'hfc, 8'h0c, 8'h0d, 8'h0c, 8'h07, 8'hf1, 8'h12, 8'h10, 8'h03, 8'h0a, 8'hf5, 8'hf1, 8'he8, 8'hff, 8'h1c, 8'h0f, 8'hf7, 8'h0a, 8'he0, 8'hef, 8'h0b, 8'hef, 8'h15, 8'hf4, 8'hfa, 8'hf5, 8'hff, 8'hf5, 8'h0c, 8'hf1, 8'h08, 8'h0c, 8'h2a, 8'h11, 8'hf0, 8'hf1, 8'hfa, 8'hf5, 8'h04, 8'he2, 8'h12, 8'h05, 8'h16, 8'hf6, 8'h0e, 8'h16, 8'h15, 8'hf4, 8'hfd, 8'h07, 8'h0f, 8'h17, 8'h04};
assign weight_matrix[81] = {8'hee, 8'h02, 8'hf4, 8'h12, 8'h0c, 8'h00, 8'hfb, 8'hf8, 8'h21, 8'h04, 8'h0e, 8'hf0, 8'h04, 8'h07, 8'h17, 8'hff, 8'hf0, 8'h0d, 8'h10, 8'hf9, 8'hea, 8'h08, 8'h07, 8'he4, 8'h00, 8'hfa, 8'hfe, 8'h0c, 8'h0d, 8'hfd, 8'hf0, 8'h17, 8'hf2, 8'hf3, 8'h04, 8'h0d, 8'hff, 8'h07, 8'h0c, 8'h02, 8'hf3, 8'hf4, 8'h0e, 8'h0b, 8'hfa, 8'h08, 8'h16, 8'hf1, 8'h03, 8'hf2, 8'h09, 8'hef, 8'h1b, 8'hf2, 8'h17, 8'h0e, 8'hfc, 8'hec, 8'h0e, 8'hf9, 8'hf4, 8'hec, 8'h15, 8'h18};
assign weight_matrix[82] = {8'h06, 8'hf5, 8'h0e, 8'hec, 8'hf1, 8'hf8, 8'hf4, 8'h0e, 8'hfd, 8'hf3, 8'hf5, 8'h13, 8'h0f, 8'h0a, 8'h0a, 8'hf8, 8'h10, 8'hf8, 8'h10, 8'h0a, 8'hf9, 8'h12, 8'h0b, 8'h08, 8'hfa, 8'h09, 8'h0f, 8'hfe, 8'h13, 8'hee, 8'h00, 8'hff, 8'h08, 8'h14, 8'hec, 8'hf0, 8'hea, 8'hf7, 8'hf7, 8'hea, 8'h0d, 8'hf5, 8'h06, 8'h00, 8'h09, 8'hf4, 8'h08, 8'hf8, 8'h06, 8'h0f, 8'hf6, 8'h10, 8'hef, 8'h07, 8'hf8, 8'hee, 8'hfd, 8'h12, 8'hff, 8'hf9, 8'hfb, 8'hfa, 8'hfd, 8'h01};
assign weight_matrix[83] = {8'hf5, 8'h12, 8'h15, 8'h13, 8'hf2, 8'h0d, 8'hf0, 8'hfb, 8'hf6, 8'hf6, 8'h0b, 8'he9, 8'hed, 8'hf0, 8'h0d, 8'h09, 8'h14, 8'h15, 8'h0e, 8'hf4, 8'hfd, 8'hfa, 8'h00, 8'h07, 8'h04, 8'h08, 8'h02, 8'h0d, 8'h0d, 8'h12, 8'h05, 8'h0c, 8'hf4, 8'h0e, 8'hf6, 8'h10, 8'h05, 8'h0d, 8'heb, 8'hfe, 8'hef, 8'h13, 8'hf9, 8'hf6, 8'h14, 8'h11, 8'h13, 8'h11, 8'h00, 8'hfc, 8'h12, 8'hfb, 8'h00, 8'h0f, 8'h00, 8'h13, 8'heb, 8'hef, 8'h09, 8'hee, 8'hee, 8'h0a, 8'h04, 8'hf4};
assign weight_matrix[84] = {8'h06, 8'hfa, 8'h04, 8'h0f, 8'h08, 8'h02, 8'h11, 8'he8, 8'hfe, 8'h0a, 8'h19, 8'h03, 8'he0, 8'h0c, 8'hea, 8'h06, 8'h0a, 8'hf9, 8'hf8, 8'hf8, 8'hfc, 8'h13, 8'h06, 8'hf9, 8'he7, 8'h13, 8'hf7, 8'h0b, 8'hf6, 8'h16, 8'hf9, 8'hf2, 8'h0a, 8'he3, 8'h03, 8'hfc, 8'he5, 8'h02, 8'h04, 8'hf3, 8'h0e, 8'h03, 8'hf9, 8'hf0, 8'h1b, 8'hf9, 8'hf5, 8'h0c, 8'hfa, 8'h03, 8'h1d, 8'he6, 8'hfa, 8'h16, 8'hfc, 8'hfc, 8'hfd, 8'h27, 8'h02, 8'hfc, 8'hec, 8'h0e, 8'h00, 8'hd8};
assign weight_matrix[85] = {8'hf7, 8'hff, 8'h10, 8'hf5, 8'hf6, 8'hf9, 8'h03, 8'h06, 8'h0b, 8'hec, 8'hee, 8'hf4, 8'hfc, 8'h07, 8'hec, 8'h00, 8'h04, 8'hfa, 8'hf4, 8'h0a, 8'hf2, 8'h16, 8'hee, 8'hf0, 8'h0d, 8'h0d, 8'h0d, 8'hfe, 8'hfc, 8'h04, 8'h02, 8'h07, 8'hf3, 8'h00, 8'hf9, 8'h0c, 8'hf3, 8'hfe, 8'h14, 8'h12, 8'h0e, 8'h01, 8'h11, 8'h02, 8'h13, 8'h11, 8'h10, 8'h10, 8'hfc, 8'hf3, 8'h10, 8'hec, 8'h06, 8'hfa, 8'heb, 8'h05, 8'h09, 8'h0c, 8'hfd, 8'h0d, 8'h09, 8'hee, 8'h15, 8'h14};
assign weight_matrix[86] = {8'h0a, 8'h0c, 8'hf1, 8'hff, 8'hed, 8'h11, 8'hfa, 8'h0a, 8'h11, 8'h08, 8'hf9, 8'h12, 8'h12, 8'hf1, 8'hed, 8'hec, 8'hf0, 8'hfe, 8'h00, 8'hff, 8'hef, 8'hed, 8'hfe, 8'hf5, 8'h01, 8'h04, 8'hea, 8'hfb, 8'hf5, 8'h0e, 8'hec, 8'hfd, 8'hf9, 8'hec, 8'heb, 8'h09, 8'h0c, 8'hfd, 8'h0f, 8'h07, 8'h03, 8'hfb, 8'h0b, 8'h07, 8'hee, 8'h04, 8'h0e, 8'hf3, 8'h13, 8'heb, 8'h13, 8'h00, 8'he9, 8'hff, 8'hf7, 8'heb, 8'he9, 8'hf0, 8'h02, 8'hf3, 8'h01, 8'hfe, 8'h03, 8'hf5};
assign weight_matrix[87] = {8'h00, 8'h04, 8'hff, 8'h0a, 8'h0a, 8'h0b, 8'hec, 8'hfb, 8'hf7, 8'h0f, 8'h05, 8'h02, 8'hfe, 8'hea, 8'hfe, 8'h05, 8'h00, 8'hf0, 8'h13, 8'hf7, 8'h09, 8'h07, 8'h0b, 8'hfc, 8'h12, 8'hfd, 8'h12, 8'h02, 8'hee, 8'hf2, 8'hfe, 8'hf1, 8'h01, 8'hf3, 8'h06, 8'heb, 8'h06, 8'hf4, 8'hf6, 8'hff, 8'hfc, 8'h11, 8'h0c, 8'hfc, 8'hfe, 8'hea, 8'h0e, 8'h09, 8'h0f, 8'h13, 8'h08, 8'hec, 8'h05, 8'h10, 8'hf7, 8'hf8, 8'h07, 8'hf3, 8'h00, 8'h14, 8'hea, 8'h0e, 8'h0d, 8'h06};
assign weight_matrix[88] = {8'h0b, 8'hfb, 8'h09, 8'h0a, 8'hef, 8'hee, 8'hea, 8'h0f, 8'h0c, 8'h13, 8'hfd, 8'h04, 8'hf4, 8'h09, 8'h0f, 8'hf3, 8'hf8, 8'hff, 8'hf6, 8'hf8, 8'hfa, 8'hf6, 8'h00, 8'hed, 8'hf8, 8'hfd, 8'hf9, 8'h07, 8'h11, 8'h00, 8'hfb, 8'hf4, 8'h18, 8'h0d, 8'hec, 8'h03, 8'hf0, 8'hea, 8'hfe, 8'hf9, 8'hfc, 8'h10, 8'h13, 8'h10, 8'h0b, 8'hf9, 8'hfe, 8'hfa, 8'hf2, 8'h13, 8'h13, 8'hef, 8'h01, 8'h07, 8'hf1, 8'h12, 8'hf7, 8'hed, 8'hff, 8'h0e, 8'hf4, 8'h05, 8'hfa, 8'hf0};
assign weight_matrix[89] = {8'he9, 8'he4, 8'h0a, 8'hea, 8'h0a, 8'h0b, 8'hed, 8'hf0, 8'h19, 8'h2a, 8'he7, 8'h10, 8'hf5, 8'h07, 8'heb, 8'h02, 8'h13, 8'hee, 8'h09, 8'hf3, 8'hec, 8'h05, 8'h07, 8'h12, 8'h0c, 8'he4, 8'h13, 8'hf6, 8'hec, 8'h1d, 8'h05, 8'h00, 8'h2a, 8'hf8, 8'h0c, 8'hea, 8'hff, 8'h02, 8'he4, 8'hf1, 8'hf3, 8'hec, 8'heb, 8'hd2, 8'h17, 8'h12, 8'hef, 8'h05, 8'hed, 8'h06, 8'h11, 8'hee, 8'hf9, 8'he0, 8'h17, 8'hf7, 8'hff, 8'h09, 8'hfe, 8'hec, 8'h09, 8'h19, 8'hf4, 8'he7};
assign weight_matrix[90] = {8'hf5, 8'hf6, 8'hf5, 8'h10, 8'hf5, 8'hf4, 8'h0e, 8'hea, 8'h03, 8'he8, 8'h03, 8'heb, 8'h10, 8'he6, 8'hf0, 8'h04, 8'hee, 8'h03, 8'h0b, 8'heb, 8'h0c, 8'hf6, 8'h03, 8'h02, 8'h0c, 8'hd5, 8'hea, 8'hf3, 8'hef, 8'hf9, 8'h10, 8'h11, 8'hf7, 8'h0a, 8'h14, 8'hfc, 8'h05, 8'hf3, 8'h08, 8'h02, 8'h0e, 8'h08, 8'h11, 8'h0c, 8'h11, 8'hed, 8'hf6, 8'hfb, 8'h01, 8'hfa, 8'hf0, 8'h19, 8'hf9, 8'h01, 8'hfd, 8'hf1, 8'h09, 8'he3, 8'h0b, 8'h0b, 8'h04, 8'he5, 8'h05, 8'h27};
assign weight_matrix[91] = {8'h00, 8'hf0, 8'h02, 8'h0c, 8'hf4, 8'h10, 8'hfd, 8'h0e, 8'h00, 8'hf0, 8'hfb, 8'hf2, 8'h04, 8'hf0, 8'hf2, 8'h0a, 8'hef, 8'hf2, 8'hf1, 8'h07, 8'h00, 8'hff, 8'hf1, 8'h05, 8'h0a, 8'hf8, 8'he8, 8'h0c, 8'h00, 8'hff, 8'h03, 8'hf1, 8'h11, 8'hfd, 8'hfe, 8'h00, 8'hea, 8'hee, 8'hf4, 8'hfa, 8'h05, 8'hfe, 8'hfe, 8'h03, 8'hee, 8'h00, 8'hfb, 8'hf9, 8'he8, 8'hf8, 8'h00, 8'hf1, 8'h01, 8'h0e, 8'h00, 8'h0c, 8'hfb, 8'hf9, 8'he3, 8'hf6, 8'hf0, 8'hf9, 8'h02, 8'h06};
assign weight_matrix[92] = {8'hed, 8'hf7, 8'h08, 8'hf9, 8'hf2, 8'hf6, 8'h0e, 8'h14, 8'h27, 8'hfc, 8'h0d, 8'he8, 8'h19, 8'h06, 8'h15, 8'h1f, 8'h04, 8'he3, 8'h0b, 8'hfd, 8'h06, 8'he5, 8'hea, 8'hef, 8'h00, 8'hee, 8'hf8, 8'hf3, 8'hf5, 8'he6, 8'hec, 8'h17, 8'hf0, 8'hfa, 8'h14, 8'hff, 8'h31, 8'h1a, 8'h1a, 8'hf1, 8'h03, 8'h04, 8'h0e, 8'h11, 8'hed, 8'hf6, 8'h05, 8'hf6, 8'hea, 8'hf7, 8'he9, 8'hf1, 8'h13, 8'hf0, 8'hf5, 8'hf8, 8'he8, 8'hde, 8'hf6, 8'hf3, 8'hf0, 8'he6, 8'h0f, 8'h24};
assign weight_matrix[93] = {8'hfd, 8'hfa, 8'h07, 8'hfe, 8'hfd, 8'hf8, 8'hf4, 8'h08, 8'h13, 8'hfe, 8'h05, 8'h14, 8'h0c, 8'hfa, 8'h04, 8'h0b, 8'heb, 8'h04, 8'hef, 8'hfc, 8'h00, 8'hf4, 8'hf9, 8'h13, 8'h09, 8'h0a, 8'h14, 8'hef, 8'h05, 8'hfd, 8'h0f, 8'h10, 8'hfc, 8'hfb, 8'hf9, 8'hfe, 8'h13, 8'h0e, 8'h05, 8'h08, 8'h0e, 8'h06, 8'hfa, 8'hf7, 8'h0a, 8'hfe, 8'h0f, 8'h16, 8'h10, 8'h11, 8'h05, 8'h06, 8'hfc, 8'hea, 8'hfa, 8'hf4, 8'hfa, 8'h11, 8'hf7, 8'hf6, 8'hf4, 8'hfd, 8'h0c, 8'hf7};
assign weight_matrix[94] = {8'h03, 8'hf1, 8'hf8, 8'h01, 8'hf8, 8'h01, 8'hf2, 8'heb, 8'h04, 8'hf0, 8'hfc, 8'hef, 8'hfc, 8'hfe, 8'hf1, 8'h0b, 8'h14, 8'hf1, 8'hf6, 8'heb, 8'h10, 8'hf8, 8'hf3, 8'h10, 8'h0f, 8'hff, 8'hf6, 8'he9, 8'hf4, 8'h11, 8'hef, 8'hf1, 8'hfe, 8'hf5, 8'hff, 8'hf0, 8'h07, 8'h10, 8'hf5, 8'hf7, 8'hea, 8'hfa, 8'hf1, 8'h08, 8'hf4, 8'hfb, 8'hf2, 8'he8, 8'h11, 8'hec, 8'h0d, 8'hfb, 8'hf1, 8'hf8, 8'hff, 8'hf9, 8'hf9, 8'hf9, 8'hff, 8'h03, 8'hfc, 8'hf6, 8'hfe, 8'h0a};
assign weight_matrix[95] = {8'h0e, 8'hfb, 8'h11, 8'hed, 8'h15, 8'h0f, 8'hd0, 8'h01, 8'hfc, 8'hf3, 8'he9, 8'h08, 8'heb, 8'h0b, 8'h17, 8'h13, 8'h00, 8'hfb, 8'h10, 8'he9, 8'h0d, 8'h03, 8'h0f, 8'h09, 8'h0e, 8'hef, 8'hf6, 8'h1a, 8'h00, 8'h15, 8'hf9, 8'hed, 8'h1a, 8'h24, 8'hee, 8'h0f, 8'h05, 8'hf3, 8'h08, 8'h0e, 8'h15, 8'hf4, 8'hfb, 8'h00, 8'h32, 8'h1c, 8'he8, 8'hfc, 8'h19, 8'hf7, 8'h14, 8'hf6, 8'h0f, 8'hf9, 8'h1a, 8'h0a, 8'hfc, 8'hf8, 8'hfb, 8'h00, 8'he8, 8'hfc, 8'hf7, 8'hf1};
assign weight_matrix[96] = {8'h02, 8'h11, 8'hea, 8'h00, 8'hfe, 8'hec, 8'h0c, 8'h05, 8'he9, 8'hf1, 8'h11, 8'h00, 8'h0b, 8'hf9, 8'h02, 8'hfa, 8'hf3, 8'hfe, 8'hea, 8'hfe, 8'hf3, 8'hf2, 8'hf9, 8'h10, 8'hfc, 8'he7, 8'h06, 8'hff, 8'hf3, 8'h19, 8'h0b, 8'h08, 8'h19, 8'he9, 8'h05, 8'hea, 8'hef, 8'h04, 8'h06, 8'hfe, 8'h15, 8'h04, 8'h0e, 8'hea, 8'h0d, 8'hf2, 8'hf6, 8'h08, 8'hea, 8'hef, 8'hfe, 8'hfd, 8'hfa, 8'h09, 8'h07, 8'hf0, 8'hff, 8'hfe, 8'hfc, 8'hf5, 8'hf6, 8'hf3, 8'h0a, 8'h11};
assign weight_matrix[97] = {8'hf8, 8'h02, 8'h0e, 8'h02, 8'h01, 8'hef, 8'hf4, 8'hf4, 8'hef, 8'hfe, 8'h0f, 8'h14, 8'h00, 8'h13, 8'h05, 8'hf3, 8'h19, 8'heb, 8'hf2, 8'h14, 8'hee, 8'h15, 8'hf1, 8'h0c, 8'h0d, 8'heb, 8'h12, 8'h14, 8'h16, 8'h13, 8'hec, 8'h11, 8'hf0, 8'hf8, 8'hf2, 8'hf8, 8'h0d, 8'hea, 8'hf1, 8'h07, 8'hf9, 8'h04, 8'h11, 8'hec, 8'hfb, 8'h00, 8'h0c, 8'h02, 8'h03, 8'hf7, 8'h01, 8'hf6, 8'h13, 8'hf4, 8'h21, 8'h0a, 8'h03, 8'heb, 8'hf7, 8'hf7, 8'h10, 8'h09, 8'hfd, 8'hef};
assign weight_matrix[98] = {8'h0a, 8'hf6, 8'hf4, 8'h0c, 8'h11, 8'hf4, 8'hf7, 8'hf2, 8'hf6, 8'hf3, 8'h07, 8'h0f, 8'hf3, 8'hfb, 8'hf7, 8'hfc, 8'h0f, 8'hf8, 8'hfc, 8'hed, 8'h11, 8'hf5, 8'h02, 8'hfe, 8'h10, 8'h14, 8'h02, 8'h0f, 8'hf9, 8'hfc, 8'h00, 8'h00, 8'hf0, 8'h10, 8'hfc, 8'heb, 8'h01, 8'hf6, 8'h01, 8'h0d, 8'h0f, 8'h12, 8'hfe, 8'hf1, 8'h16, 8'hf6, 8'h0e, 8'h0c, 8'h03, 8'h03, 8'h03, 8'hf4, 8'h0b, 8'hf2, 8'h09, 8'h0d, 8'hfe, 8'h10, 8'h00, 8'h13, 8'hf7, 8'hfc, 8'hf8, 8'hee};
assign weight_matrix[99] = {8'h06, 8'hf2, 8'h12, 8'h16, 8'hf6, 8'hec, 8'h09, 8'h0f, 8'h00, 8'h08, 8'hff, 8'h11, 8'hf2, 8'hed, 8'h04, 8'hf2, 8'h04, 8'h11, 8'hf6, 8'hf2, 8'hfc, 8'hf1, 8'hf4, 8'h13, 8'hfc, 8'h10, 8'hfa, 8'h0d, 8'h0f, 8'h09, 8'hf3, 8'h01, 8'hfa, 8'hfc, 8'hf7, 8'h15, 8'h0a, 8'hfa, 8'h00, 8'h0b, 8'h06, 8'hf0, 8'h13, 8'h00, 8'hf5, 8'hf0, 8'h00, 8'hf7, 8'hf2, 8'heb, 8'hff, 8'h07, 8'hea, 8'hf9, 8'hf7, 8'hf5, 8'h0e, 8'h0c, 8'hf1, 8'hf7, 8'h09, 8'h0c, 8'h0c, 8'hfe};
assign weight_matrix[100] = {8'hce, 8'h14, 8'h00, 8'heb, 8'hfd, 8'hff, 8'he9, 8'heb, 8'h03, 8'h06, 8'hf7, 8'hec, 8'hef, 8'hfd, 8'h05, 8'hf3, 8'h11, 8'h10, 8'hef, 8'hff, 8'hfe, 8'hee, 8'hfe, 8'h15, 8'hf2, 8'h13, 8'h09, 8'hf6, 8'hf3, 8'h08, 8'h0b, 8'hea, 8'h16, 8'he5, 8'hf8, 8'h0a, 8'hea, 8'hf5, 8'hfe, 8'h10, 8'h00, 8'hfc, 8'h0c, 8'heb, 8'hf8, 8'h03, 8'he6, 8'hf7, 8'h0b, 8'hfb, 8'hfb, 8'hf4, 8'h0d, 8'h02, 8'h15, 8'hfd, 8'hef, 8'h23, 8'h06, 8'hfc, 8'he5, 8'h24, 8'hd3, 8'hcb};
assign weight_matrix[101] = {8'hf4, 8'hf6, 8'hee, 8'hfe, 8'hea, 8'hec, 8'hfb, 8'h11, 8'h04, 8'hf8, 8'hfa, 8'h00, 8'hf3, 8'hfc, 8'h00, 8'he7, 8'hf1, 8'hed, 8'h0a, 8'hfe, 8'hea, 8'hef, 8'hfb, 8'h0e, 8'h01, 8'h02, 8'hf3, 8'hf4, 8'h0b, 8'h0a, 8'hea, 8'hed, 8'h09, 8'hf2, 8'hfe, 8'h0a, 8'he9, 8'hfb, 8'h06, 8'he7, 8'hf6, 8'hea, 8'h10, 8'hf9, 8'hf8, 8'h0f, 8'hf3, 8'h08, 8'h0d, 8'h01, 8'hee, 8'h0e, 8'h11, 8'h0b, 8'hf7, 8'hef, 8'h0c, 8'hf3, 8'hee, 8'hef, 8'hef, 8'h09, 8'h12, 8'h00};
assign weight_matrix[102] = {8'hf0, 8'hf2, 8'h0c, 8'hfa, 8'hea, 8'hf4, 8'h01, 8'h11, 8'hee, 8'hf3, 8'hed, 8'h06, 8'h08, 8'h03, 8'hee, 8'hfb, 8'hec, 8'h09, 8'h0a, 8'h0d, 8'h09, 8'h09, 8'hfb, 8'hec, 8'hfa, 8'heb, 8'hec, 8'hf3, 8'hf5, 8'h12, 8'hf1, 8'hed, 8'hfc, 8'hf0, 8'hf6, 8'h05, 8'h0f, 8'h09, 8'hef, 8'h01, 8'h0e, 8'h07, 8'h0e, 8'h0e, 8'h16, 8'hff, 8'hf4, 8'hf8, 8'hf4, 8'h13, 8'hf7, 8'h10, 8'h11, 8'hf0, 8'h02, 8'h16, 8'hf9, 8'h0d, 8'hef, 8'hff, 8'h12, 8'hed, 8'h0f, 8'h00};
assign weight_matrix[103] = {8'h15, 8'hf4, 8'h16, 8'hfc, 8'hf6, 8'hfa, 8'hf4, 8'hfc, 8'h12, 8'hfb, 8'hf7, 8'hfd, 8'heb, 8'h11, 8'hfc, 8'h00, 8'h0a, 8'hfc, 8'h0d, 8'hf6, 8'h09, 8'h13, 8'hf6, 8'hed, 8'h15, 8'h15, 8'h0d, 8'h15, 8'hf2, 8'h02, 8'h07, 8'h0f, 8'hee, 8'hf8, 8'hf0, 8'h06, 8'h10, 8'h12, 8'h00, 8'hf3, 8'hed, 8'hfb, 8'h10, 8'h05, 8'hf6, 8'hf1, 8'hff, 8'h08, 8'h05, 8'h10, 8'hf2, 8'hec, 8'h13, 8'hed, 8'h03, 8'h15, 8'h05, 8'h0e, 8'hfd, 8'hea, 8'h02, 8'hf2, 8'h16, 8'h15};
assign weight_matrix[104] = {8'hf9, 8'h0f, 8'hf8, 8'h00, 8'hea, 8'hf8, 8'h19, 8'hf6, 8'h07, 8'hf9, 8'hf3, 8'hfd, 8'hfe, 8'h0f, 8'h0b, 8'he9, 8'hf6, 8'hee, 8'h02, 8'hff, 8'h0c, 8'hf6, 8'h01, 8'hef, 8'hfe, 8'hfd, 8'hf0, 8'h07, 8'h09, 8'hf5, 8'h0c, 8'h07, 8'h04, 8'hf4, 8'hee, 8'hf6, 8'hec, 8'h05, 8'h00, 8'hf2, 8'h0e, 8'h0c, 8'h05, 8'hf8, 8'hf3, 8'heb, 8'h06, 8'he9, 8'he9, 8'h14, 8'hf4, 8'h10, 8'h08, 8'hef, 8'hfb, 8'h02, 8'hf8, 8'h13, 8'h0e, 8'hf7, 8'h07, 8'h04, 8'hfc, 8'hf1};
assign weight_matrix[105] = {8'h03, 8'h13, 8'h09, 8'hf2, 8'hfc, 8'he9, 8'h02, 8'h0b, 8'h0c, 8'hf2, 8'hf2, 8'hed, 8'h0a, 8'h11, 8'he8, 8'h0f, 8'hfa, 8'h0a, 8'hf7, 8'h08, 8'hf1, 8'h11, 8'hff, 8'h00, 8'hf4, 8'hea, 8'hf0, 8'h11, 8'h00, 8'h0f, 8'hf8, 8'hf4, 8'hf4, 8'hf9, 8'h0f, 8'h05, 8'h13, 8'h03, 8'hf6, 8'hfe, 8'h0d, 8'h0e, 8'h07, 8'hf1, 8'h0f, 8'h09, 8'hf0, 8'hf3, 8'hfa, 8'h0a, 8'h14, 8'hf2, 8'hf3, 8'h11, 8'hf8, 8'h02, 8'h08, 8'hee, 8'he5, 8'hf1, 8'h0f, 8'hee, 8'h0a, 8'hf2};
assign weight_matrix[106] = {8'h08, 8'h06, 8'h09, 8'h07, 8'hf1, 8'h04, 8'hef, 8'h11, 8'hfd, 8'h13, 8'h13, 8'hfa, 8'hfb, 8'hf2, 8'h0d, 8'hea, 8'h08, 8'h11, 8'h0c, 8'h0d, 8'heb, 8'h03, 8'h11, 8'hfb, 8'hf0, 8'h0a, 8'h0b, 8'h09, 8'h00, 8'hf7, 8'h03, 8'hf9, 8'h0e, 8'h0d, 8'h0b, 8'h06, 8'heb, 8'hf6, 8'hfa, 8'hea, 8'h02, 8'hef, 8'hec, 8'h07, 8'h08, 8'hef, 8'h05, 8'hf8, 8'hfb, 8'hfb, 8'hf9, 8'hf0, 8'h08, 8'h09, 8'h0a, 8'hfa, 8'hfb, 8'h08, 8'h15, 8'he9, 8'hfc, 8'h0c, 8'h04, 8'hf9};
assign weight_matrix[107] = {8'h00, 8'h02, 8'hf6, 8'hff, 8'h12, 8'hf3, 8'h02, 8'h06, 8'h0f, 8'hfc, 8'h05, 8'hef, 8'hf9, 8'h0f, 8'he9, 8'hed, 8'hf2, 8'h08, 8'h07, 8'hfc, 8'hfb, 8'h03, 8'hfe, 8'h1d, 8'h0d, 8'h09, 8'h12, 8'h04, 8'h0f, 8'h1c, 8'h05, 8'hf7, 8'h17, 8'h14, 8'h07, 8'hf2, 8'h02, 8'hee, 8'he9, 8'hfd, 8'hff, 8'hf5, 8'hf8, 8'he4, 8'h03, 8'hff, 8'h0e, 8'h04, 8'hf0, 8'h08, 8'h17, 8'hf1, 8'hf9, 8'he7, 8'h10, 8'hec, 8'h04, 8'h17, 8'h10, 8'h02, 8'h05, 8'h1a, 8'hed, 8'h02};
assign weight_matrix[108] = {8'hf6, 8'heb, 8'hfb, 8'hf7, 8'h0e, 8'heb, 8'h0e, 8'h12, 8'hea, 8'h00, 8'hfe, 8'h13, 8'h0e, 8'hef, 8'hf6, 8'h08, 8'h00, 8'h11, 8'h13, 8'hf7, 8'hf5, 8'hf2, 8'hfb, 8'he9, 8'h06, 8'hf6, 8'hfa, 8'hed, 8'h06, 8'hf6, 8'h10, 8'hfb, 8'hfa, 8'h08, 8'h00, 8'hf1, 8'h0f, 8'hf8, 8'he7, 8'hf3, 8'h0a, 8'h0a, 8'hed, 8'hf3, 8'h04, 8'hff, 8'h05, 8'h04, 8'h0c, 8'heb, 8'h13, 8'hfa, 8'heb, 8'hfb, 8'h09, 8'he7, 8'h0e, 8'hed, 8'hfe, 8'hfa, 8'h06, 8'hfe, 8'h03, 8'hf6};
assign weight_matrix[109] = {8'hf5, 8'hf4, 8'hf5, 8'h10, 8'hfb, 8'h16, 8'hff, 8'hf5, 8'h0b, 8'hf7, 8'hff, 8'hfb, 8'heb, 8'h0d, 8'hf3, 8'hf9, 8'h11, 8'hfc, 8'h01, 8'h12, 8'h13, 8'h12, 8'h11, 8'hf8, 8'hfa, 8'hef, 8'h03, 8'hfc, 8'h10, 8'h13, 8'h08, 8'h08, 8'hf4, 8'hee, 8'h11, 8'h16, 8'hec, 8'h06, 8'hfa, 8'h0b, 8'hf7, 8'h02, 8'hf9, 8'h0b, 8'hed, 8'hff, 8'h15, 8'hf9, 8'h09, 8'hfe, 8'h09, 8'h12, 8'hf3, 8'hf3, 8'h0c, 8'hf1, 8'hfe, 8'h03, 8'h11, 8'hf5, 8'h05, 8'hf1, 8'h0c, 8'h13};
assign weight_matrix[110] = {8'h15, 8'hfc, 8'hf8, 8'hf1, 8'h03, 8'h11, 8'h0f, 8'h04, 8'h04, 8'h18, 8'he7, 8'hee, 8'hf6, 8'hf5, 8'hf4, 8'heb, 8'hf9, 8'h06, 8'h0a, 8'he6, 8'hf4, 8'h05, 8'hfa, 8'hff, 8'h01, 8'hd4, 8'h06, 8'hec, 8'hf0, 8'h07, 8'hf1, 8'h18, 8'h0e, 8'h0e, 8'hfd, 8'h08, 8'hec, 8'hec, 8'hf2, 8'h13, 8'hf3, 8'h05, 8'he7, 8'hfa, 8'h01, 8'hf3, 8'h07, 8'h07, 8'hf2, 8'h14, 8'h10, 8'hfe, 8'hfe, 8'he6, 8'h10, 8'h00, 8'h0e, 8'hde, 8'h12, 8'h02, 8'hf0, 8'hec, 8'h0f, 8'h1d};
assign weight_matrix[111] = {8'h0b, 8'h04, 8'hfc, 8'h06, 8'hf8, 8'h0c, 8'hea, 8'hf6, 8'hf2, 8'hf0, 8'hf7, 8'h0d, 8'hf6, 8'heb, 8'hea, 8'h04, 8'h10, 8'h00, 8'hf1, 8'h09, 8'hef, 8'hf5, 8'hfe, 8'h01, 8'h07, 8'h09, 8'hfc, 8'h01, 8'h12, 8'hf1, 8'h02, 8'h08, 8'h01, 8'hee, 8'h0e, 8'h06, 8'hf2, 8'hf7, 8'hf1, 8'hf2, 8'hf0, 8'hff, 8'h05, 8'hfa, 8'hfc, 8'hf0, 8'hf1, 8'hf2, 8'hf5, 8'hfe, 8'hf6, 8'h09, 8'h12, 8'hf3, 8'h04, 8'hef, 8'h0f, 8'h0f, 8'hed, 8'hfc, 8'h12, 8'h13, 8'h04, 8'h0d};
assign weight_matrix[112] = {8'hfa, 8'h03, 8'hef, 8'hf8, 8'hff, 8'h02, 8'h02, 8'hf8, 8'h09, 8'hed, 8'hee, 8'h10, 8'h13, 8'hfa, 8'h05, 8'h01, 8'h12, 8'hfb, 8'hf8, 8'hf6, 8'h10, 8'hf3, 8'hf5, 8'hec, 8'hf8, 8'h02, 8'h12, 8'hf1, 8'h11, 8'h08, 8'hf6, 8'hff, 8'hf4, 8'h12, 8'hec, 8'hef, 8'h0d, 8'hff, 8'hfa, 8'h0c, 8'hf9, 8'h03, 8'h13, 8'hf7, 8'h14, 8'h13, 8'hff, 8'h10, 8'hf7, 8'hef, 8'hf1, 8'hf9, 8'h0a, 8'hee, 8'hea, 8'hfd, 8'h0c, 8'h0c, 8'h0b, 8'h07, 8'hf4, 8'hec, 8'h03, 8'hf5};
assign weight_matrix[113] = {8'h04, 8'h0e, 8'h10, 8'h01, 8'h07, 8'h05, 8'he6, 8'hea, 8'hf6, 8'h0c, 8'hf4, 8'hff, 8'h0d, 8'h03, 8'hec, 8'hea, 8'h03, 8'hec, 8'hfe, 8'hff, 8'hf7, 8'h08, 8'hfb, 8'h05, 8'hfb, 8'h0c, 8'h03, 8'h08, 8'hf6, 8'h14, 8'h0c, 8'hfb, 8'hf7, 8'h03, 8'heb, 8'h11, 8'hfa, 8'h01, 8'hf5, 8'h00, 8'h0e, 8'hf3, 8'hf3, 8'h0d, 8'hf6, 8'hfd, 8'hed, 8'h08, 8'hfe, 8'h0a, 8'hfa, 8'h04, 8'he8, 8'hef, 8'h0f, 8'h04, 8'h02, 8'hf3, 8'hfa, 8'hfc, 8'hf9, 8'h05, 8'hfb, 8'hf9};
assign weight_matrix[114] = {8'hfc, 8'hf9, 8'hfc, 8'hf8, 8'h09, 8'hf8, 8'hf9, 8'h10, 8'hf5, 8'h05, 8'h14, 8'h13, 8'hfb, 8'hfb, 8'h02, 8'he8, 8'h08, 8'hfe, 8'hf0, 8'h04, 8'h03, 8'he8, 8'hea, 8'h00, 8'hfa, 8'hfb, 8'hf7, 8'hf6, 8'hee, 8'h08, 8'h06, 8'hf1, 8'hf4, 8'hfe, 8'h03, 8'hf9, 8'hfc, 8'h00, 8'h0a, 8'h03, 8'heb, 8'h06, 8'h04, 8'h06, 8'h09, 8'h09, 8'hfc, 8'hec, 8'hf6, 8'hf8, 8'h09, 8'h0b, 8'h11, 8'h08, 8'h07, 8'h08, 8'h00, 8'h0d, 8'h0f, 8'he9, 8'h10, 8'hf1, 8'hf5, 8'h00};
assign weight_matrix[115] = {8'he8, 8'hf9, 8'h0d, 8'h02, 8'h16, 8'hf5, 8'h00, 8'hff, 8'hee, 8'h0b, 8'h06, 8'hea, 8'h0e, 8'h05, 8'hf3, 8'h08, 8'h10, 8'hfd, 8'hef, 8'h0f, 8'h10, 8'hea, 8'h0c, 8'h0d, 8'h10, 8'h01, 8'hfb, 8'heb, 8'h06, 8'h10, 8'h11, 8'hfc, 8'h1d, 8'h01, 8'h06, 8'h0e, 8'hf9, 8'hfb, 8'hec, 8'hf0, 8'hf7, 8'h1d, 8'hfa, 8'hec, 8'h03, 8'h08, 8'hfa, 8'hf8, 8'h01, 8'hfa, 8'h06, 8'hf8, 8'h16, 8'h0f, 8'h0d, 8'hee, 8'h0a, 8'h17, 8'h15, 8'hfb, 8'hfe, 8'h16, 8'hee, 8'hef};
assign weight_matrix[116] = {8'h0a, 8'hfa, 8'hf6, 8'hfe, 8'h02, 8'h0c, 8'hf6, 8'he9, 8'hed, 8'hf2, 8'hed, 8'hf5, 8'h02, 8'hfc, 8'hf1, 8'hff, 8'hf4, 8'h09, 8'h0c, 8'hf5, 8'hfa, 8'h0e, 8'hfa, 8'h03, 8'hee, 8'h08, 8'hf4, 8'hf6, 8'h02, 8'hf7, 8'h09, 8'h17, 8'hf9, 8'hee, 8'h03, 8'h0b, 8'h08, 8'hf0, 8'hed, 8'hee, 8'hf8, 8'h01, 8'hf0, 8'h12, 8'hf6, 8'h05, 8'hee, 8'h08, 8'h01, 8'h00, 8'hf4, 8'hf1, 8'hf7, 8'hec, 8'h00, 8'h07, 8'hfd, 8'h0d, 8'heb, 8'hee, 8'hf3, 8'hf0, 8'hf4, 8'hfb};
assign weight_matrix[117] = {8'he4, 8'h13, 8'hdd, 8'h06, 8'hee, 8'hf7, 8'he7, 8'h04, 8'h13, 8'hec, 8'hfe, 8'hfa, 8'hf3, 8'hf6, 8'hf4, 8'h05, 8'hf0, 8'hf5, 8'hf4, 8'hec, 8'h0b, 8'hfc, 8'h06, 8'hf8, 8'hec, 8'hfd, 8'h0a, 8'hf5, 8'hf2, 8'h09, 8'hf5, 8'h12, 8'he3, 8'hff, 8'hf3, 8'h01, 8'h11, 8'h04, 8'h0c, 8'h0d, 8'h02, 8'hec, 8'hf2, 8'h35, 8'hfe, 8'hff, 8'h04, 8'h10, 8'hed, 8'h04, 8'hec, 8'h02, 8'hea, 8'hff, 8'he0, 8'h0b, 8'hee, 8'hfe, 8'h06, 8'h07, 8'hf8, 8'h02, 8'h04, 8'h02};
assign weight_matrix[118] = {8'h08, 8'hfa, 8'hfc, 8'h01, 8'hf3, 8'h0c, 8'h11, 8'heb, 8'hff, 8'hfc, 8'h16, 8'hf4, 8'h07, 8'h12, 8'h00, 8'h00, 8'h15, 8'hee, 8'hf0, 8'h0e, 8'hef, 8'hfd, 8'h08, 8'hfe, 8'hfe, 8'heb, 8'h16, 8'heb, 8'h0f, 8'h01, 8'hfd, 8'h10, 8'hf0, 8'h11, 8'hf8, 8'h12, 8'h06, 8'h12, 8'h12, 8'h14, 8'h05, 8'hfb, 8'hf4, 8'hed, 8'h11, 8'h05, 8'hfc, 8'heb, 8'h05, 8'hec, 8'h15, 8'hed, 8'hfd, 8'hff, 8'h05, 8'h08, 8'h01, 8'hed, 8'hec, 8'hf8, 8'h0a, 8'hf7, 8'hf1, 8'hff};
assign weight_matrix[119] = {8'h0f, 8'hf2, 8'heb, 8'hf0, 8'hef, 8'hf8, 8'hed, 8'hf9, 8'hfc, 8'h09, 8'hff, 8'hfa, 8'hf8, 8'hef, 8'h04, 8'h0e, 8'hfe, 8'hf5, 8'h05, 8'hf3, 8'h00, 8'hf2, 8'hed, 8'h0a, 8'hf3, 8'hfd, 8'h11, 8'hee, 8'h14, 8'h05, 8'h13, 8'h0f, 8'hff, 8'h0e, 8'h0f, 8'hfc, 8'h0c, 8'hf1, 8'h03, 8'hea, 8'h0f, 8'h03, 8'h05, 8'h01, 8'h04, 8'h00, 8'h07, 8'hf2, 8'h12, 8'h0a, 8'hf2, 8'h01, 8'h07, 8'hfa, 8'h01, 8'h0b, 8'h11, 8'h04, 8'hfe, 8'hf5, 8'h07, 8'h0b, 8'h00, 8'h0b};
assign weight_matrix[120] = {8'h04, 8'h08, 8'hf1, 8'h02, 8'hf1, 8'h00, 8'hf4, 8'h02, 8'hef, 8'h0c, 8'hfb, 8'hea, 8'h02, 8'hfa, 8'hf7, 8'h12, 8'h0d, 8'hf0, 8'hf7, 8'heb, 8'h0e, 8'hff, 8'hfa, 8'hfc, 8'hf0, 8'h03, 8'hf1, 8'hf8, 8'hec, 8'hfe, 8'h06, 8'h12, 8'h0e, 8'hf1, 8'hf5, 8'h05, 8'hfe, 8'h08, 8'hf0, 8'h03, 8'he9, 8'h01, 8'hed, 8'h05, 8'hfc, 8'h0e, 8'h01, 8'h0b, 8'h11, 8'h00, 8'hfc, 8'hf3, 8'h12, 8'hf3, 8'hfc, 8'hf7, 8'h07, 8'h05, 8'h0a, 8'h04, 8'hed, 8'hf9, 8'h12, 8'hf8};
assign weight_matrix[121] = {8'h03, 8'h0b, 8'h02, 8'h0f, 8'hef, 8'hfd, 8'h07, 8'hff, 8'hfb, 8'hed, 8'hf1, 8'hf0, 8'hed, 8'h0c, 8'h00, 8'heb, 8'hec, 8'h13, 8'he9, 8'heb, 8'hfb, 8'h0e, 8'hef, 8'hf8, 8'hfd, 8'hfa, 8'h09, 8'hf7, 8'h08, 8'hf9, 8'h12, 8'h08, 8'hee, 8'h0c, 8'h0d, 8'h10, 8'he8, 8'hf3, 8'hf8, 8'hed, 8'hfe, 8'hed, 8'hfa, 8'hf7, 8'hf2, 8'h00, 8'h12, 8'h0b, 8'hf0, 8'hec, 8'h01, 8'hf6, 8'hf6, 8'h11, 8'hf1, 8'h0c, 8'hfe, 8'h00, 8'hff, 8'hfe, 8'he9, 8'h14, 8'hf1, 8'hf0};
assign weight_matrix[122] = {8'hf0, 8'h18, 8'hf2, 8'h02, 8'h07, 8'hf4, 8'h00, 8'hea, 8'hff, 8'hf5, 8'hf6, 8'h03, 8'hf6, 8'h06, 8'hee, 8'hfa, 8'h0a, 8'hf5, 8'he8, 8'he8, 8'hf6, 8'h05, 8'hf3, 8'h0b, 8'h06, 8'h20, 8'hf0, 8'hfc, 8'hff, 8'hec, 8'h0a, 8'hfc, 8'hfc, 8'h0b, 8'hea, 8'hfd, 8'hee, 8'h13, 8'hf1, 8'h0b, 8'h0c, 8'h00, 8'hfe, 8'h10, 8'h0e, 8'hfd, 8'h0d, 8'h00, 8'heb, 8'h02, 8'hff, 8'h12, 8'hec, 8'h03, 8'hfd, 8'hec, 8'hf3, 8'h04, 8'hfe, 8'h0f, 8'h07, 8'hf7, 8'heb, 8'h08};
assign weight_matrix[123] = {8'h06, 8'hf9, 8'h0b, 8'hf0, 8'h00, 8'h10, 8'hed, 8'he8, 8'h02, 8'hec, 8'hfd, 8'hf8, 8'hf2, 8'h00, 8'hfa, 8'hfc, 8'hf0, 8'h06, 8'hf8, 8'hfb, 8'hfe, 8'h0d, 8'h11, 8'hea, 8'hfb, 8'h0a, 8'h04, 8'hf3, 8'heb, 8'hf0, 8'hed, 8'h05, 8'h13, 8'hf4, 8'hf7, 8'he7, 8'hfb, 8'h0e, 8'h07, 8'hf3, 8'hea, 8'h02, 8'h14, 8'h06, 8'hfe, 8'h04, 8'hf1, 8'he8, 8'hfc, 8'hf5, 8'h0a, 8'hff, 8'h0e, 8'h0b, 8'hfe, 8'h0e, 8'hfd, 8'h0d, 8'h1d, 8'h05, 8'hf9, 8'h13, 8'hef, 8'hf8};
assign weight_matrix[124] = {8'hf7, 8'h08, 8'h0a, 8'hed, 8'hee, 8'h00, 8'h03, 8'hec, 8'h14, 8'hfe, 8'hee, 8'hf4, 8'h0d, 8'hec, 8'h14, 8'h12, 8'h0d, 8'hf7, 8'hff, 8'hf4, 8'hf4, 8'h0c, 8'hea, 8'hf4, 8'h09, 8'h15, 8'h12, 8'h09, 8'h05, 8'h16, 8'h0f, 8'h01, 8'h0d, 8'hfc, 8'h11, 8'hed, 8'hf8, 8'h11, 8'h01, 8'hed, 8'heb, 8'h15, 8'heb, 8'hea, 8'hf9, 8'hfd, 8'heb, 8'hec, 8'hef, 8'h0e, 8'hf9, 8'hfe, 8'hf8, 8'hea, 8'hec, 8'h09, 8'hef, 8'h13, 8'hf7, 8'h09, 8'hed, 8'h11, 8'hf9, 8'hf8};
assign weight_matrix[125] = {8'h09, 8'h0c, 8'hf3, 8'hf7, 8'h06, 8'hff, 8'hf2, 8'h0c, 8'h0c, 8'h16, 8'hf7, 8'h15, 8'hff, 8'h02, 8'hf0, 8'h0b, 8'h14, 8'h01, 8'hec, 8'h11, 8'hfe, 8'hfd, 8'h16, 8'hea, 8'h08, 8'hf3, 8'hfa, 8'h08, 8'h08, 8'h10, 8'h05, 8'h03, 8'hed, 8'h12, 8'hf4, 8'h16, 8'h09, 8'h14, 8'hef, 8'h10, 8'hff, 8'h12, 8'hf8, 8'h05, 8'h15, 8'h01, 8'h14, 8'h11, 8'h01, 8'hf9, 8'hea, 8'h16, 8'hf3, 8'h0f, 8'hea, 8'h06, 8'hf5, 8'hf9, 8'h0b, 8'h01, 8'hee, 8'heb, 8'hf1, 8'h01};
assign weight_matrix[126] = {8'hfb, 8'h07, 8'h06, 8'h12, 8'h0b, 8'h16, 8'hf1, 8'h01, 8'h15, 8'hf2, 8'h07, 8'h15, 8'hff, 8'hf7, 8'h12, 8'hf8, 8'h06, 8'hf7, 8'hfe, 8'hf3, 8'hfb, 8'h09, 8'h09, 8'hf6, 8'hfd, 8'h0b, 8'hf5, 8'hf2, 8'hfc, 8'hfb, 8'hea, 8'hef, 8'hee, 8'h0f, 8'h13, 8'h0d, 8'h01, 8'h11, 8'hfc, 8'h06, 8'h04, 8'h00, 8'hf1, 8'hed, 8'hfc, 8'h12, 8'hff, 8'h0b, 8'h0f, 8'hea, 8'h11, 8'hfb, 8'h01, 8'heb, 8'hf6, 8'h0e, 8'hf1, 8'h15, 8'h0b, 8'h0d, 8'h06, 8'h10, 8'hfa, 8'hfe};
assign weight_matrix[127] = {8'h09, 8'h0e, 8'h0e, 8'h1b, 8'h13, 8'h0c, 8'h01, 8'hfd, 8'hdc, 8'h1f, 8'h06, 8'h03, 8'hed, 8'hfd, 8'h11, 8'hf2, 8'h24, 8'h07, 8'hf6, 8'h04, 8'hfc, 8'hfc, 8'h26, 8'h08, 8'h06, 8'he1, 8'he8, 8'hfc, 8'h03, 8'h14, 8'hfc, 8'hdc, 8'h35, 8'h05, 8'hfe, 8'h09, 8'hf1, 8'hee, 8'h05, 8'h0f, 8'h0c, 8'h17, 8'hf1, 8'hf8, 8'h18, 8'hed, 8'hf6, 8'hf8, 8'hee, 8'hf5, 8'h1d, 8'he2, 8'hf9, 8'hf7, 8'h0e, 8'he6, 8'hf7, 8'h0a, 8'h0c, 8'h0b, 8'h10, 8'hf6, 8'hfd, 8'hdc};

assign bias_vector = {8'h04, 8'hfe, 8'hf9, 8'hfc, 8'h00, 8'hfd, 8'h00, 8'hfc, 8'hfe, 8'hef, 8'h01, 8'h00, 8'h05, 8'hf9, 8'hf9, 8'hfe, 8'hfa, 8'hf6, 8'h08, 8'hf8, 8'hf8, 8'hfa, 8'hf5, 8'hf2, 8'hfa, 8'hf7, 8'hf9, 8'hf9, 8'h02, 8'hf3, 8'hfc, 8'h0f, 8'he7, 8'hfe, 8'hfe, 8'hfb, 8'hfd, 8'hf6, 8'hfc, 8'hf7, 8'hf8, 8'hfd, 8'hfb, 8'h14, 8'hfa, 8'hf7, 8'hfc, 8'hfb, 8'hf8, 8'hfc, 8'hf8, 8'h0b, 8'hfa, 8'hfe, 8'hef, 8'hfc, 8'hfc, 8'hf0, 8'h02, 8'hf4, 8'hfe, 8'hf4, 8'h12, 8'h15};

    
    always_ff @(posedge clk) begin
        if(rst) begin
            for (k = 0; k < OUT_SIZE_2; k++) 
            output_vector[k] <= '0;
            i <= '0;
        end else begin
            for (k = 0; k < OUT_SIZE_2; k++)
            output_vector[k] <= output_vector_nxt[k];
            i <= i_nxt;
    end
    end
    

    always_comb begin
        if (i < IN_SIZE_2) begin
            i_nxt = i + 1;
            for (j = 0; j < OUT_SIZE_2; j++) 
            output_vector_nxt[j] = output_vector[j] +  bias_vector[j] + input_vector[i] * weight_matrix[i][j];
        end else begin
            i_nxt = i;
            for (j = 0; j < OUT_SIZE_2; j++) begin
                if (output_vector[j] < 0) 
                    output_vector_nxt [j] = 0;
                else
                    output_vector_nxt [j] = output_vector [j];
            end
        end

        end
endmodule
