//tbd
module wrapper();




    
endmodule