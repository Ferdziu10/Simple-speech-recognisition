`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/24/2019 01:18:52 AM
// Design Name: 
// Module Name: dB_LUT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module dB_LUT(
    input [31:0] in,
    output [15:0] out,
    input on
    );
    
    logic [15:0] _out;
    
    assign out = _out;
    
    always_comb begin
        if(on) begin
            casex(in)
                32'b00000000000000000000000000000000: _out=0;
            
                32'b00000000000000000000000000000001: _out=0;              //1
            
                32'b00000000000000000000000000000010: _out=6;              //2
                
                32'b00000000000000000000000000000011: _out=10;              //3
                
                32'b00000000000000000000000000000100: _out=12;              //4
                
                32'b00000000000000000000000000000101: _out=14;              //5
                
                32'b00000000000000000000000000000110: _out=16;              //6
                
                32'b00000000000000000000000000000111: _out=17;              //7
                
                32'b00000000000000000000000000001000: _out=18;              //8
                
                32'b00000000000000000000000000001001: _out=19;              //9
                
                32'b00000000000000000000000000001010: _out=20;              //10
                
                32'b00000000000000000000000000001011: _out=21;              //11
                
                32'b0000000000000000000000000000110x: _out=22;              //12-13
                
                32'b00000000000000000000000000001110: _out=23;              //14
                
                32'b00000000000000000000000000001111: _out=24;              //15
                32'b00000000000000000000000000010000: _out=24;              //16
                
                32'b00000000000000000000000000010001: _out=25;              //17
                32'b00000000000000000000000000010010: _out=25;              //18
                
                32'b00000000000000000000000000010011: _out=26;              //19
                32'b0000000000000000000000000001010x: _out=26;              //20-21
                
                32'b0000000000000000000000000001011x: _out=27;              //22-23
                
                32'b0000000000000000000000000001100x: _out=28;              //24-25
                32'b00000000000000000000000000011010: _out=28;              //26
                
                32'b00000000000000000000000000011011: _out=29;              //27
                32'b0000000000000000000000000001110x: _out=29;              //28-29
                
                32'b0000000000000000000000000001111x: _out=30;              //30-31
                32'b0000000000000000000000000010000x: _out=30;              //32-33
                
                32'b0000000000000000000000000010001x: _out=31;              //34-35
                32'b0000000000000000000000000010010x: _out=31;              //36-37
                
                32'b0000000000000000000000000010011x: _out=32;              //38-39
                32'b0000000000000000000000000010100x: _out=32;              //40-41
                32'b00000000000000000000000000101010: _out=32;              //42
                
                32'b00000000000000000000000000101011: _out=33;              //43
                32'b000000000000000000000000001011xx: _out=33;              //44-47
                
                32'b000000000000000000000000001100xx: _out=34;              //48-51
                32'b0000000000000000000000000011010x: _out=34;              //52-53
                
                32'b0000000000000000000000000011011x: _out=35;              //54-55
                32'b000000000000000000000000001110xx: _out=35;              //56-59
                
                32'b000000000000000000000000001111xx: _out=36;              //60-63
                32'b0000000000000000000000000100000x: _out=36;              //64-65
                32'b00000000000000000000000001000010: _out=36;              //66
                
                32'b00000000000000000000000001000011: _out=37;              //67
                32'b000000000000000000000000010001xx: _out=37;              //68-71
                32'b0000000000000000000000000100100x: _out=37;              //72-73
                32'b00000000000000000000000001001010: _out=37;              //74
                
                32'b00000000000000000000000001001011: _out=38;              //75
                32'b100000000000000000000000000011xx: _out=38;              //76-79
                32'b000000000000000000000000010100xx: _out=38;              //80-83
                32'b00000000000000000000000001010100: _out=38;              //84
                
                32'b00000000000000000000000001010101: _out=39;              //85
                32'b0000000000000000000000000101011x: _out=39;              //86-87
                32'b000000000000000000000000010110xx: _out=39;              //88-91
                32'b0000000000000000000000000101110x: _out=39;              //92-93
                32'b00000000000000000000000001011110: _out=39;              //94
                
                32'b00000000000000000000000001011111: _out=40;              //95
                32'b00000000000000000000000001100xxx: _out=40;              //96-103
                32'b0000000000000000000000000110100x: _out=40;              //104-105
                
                32'b0000000000000000000000000110101x: _out=41;              //106-107
                32'b000000000000000000000000011011xx: _out=41;              //108-111
                32'b000000000000000000000000011100xx: _out=41;              //112-115
                32'b0000000000000000000000000111010x: _out=41;              //116-117
                32'b00000000000000000000000001110110: _out=41;              //118
                
                32'b00000000000000000000000001110111: _out=42;              //119
                32'b00000000000000000000000001111xxx: _out=42;              //120-127
                32'b000000000000000000000000100000xx: _out=42;              //128-131
                32'b0000000000000000000000001000010x: _out=42;              //132-133
                
                32'b0000000000000000000000001000011x: _out=43;              //134-135
                32'b00000000000000000000000010001xxx: _out=43;              //136-143
                32'b000000000000000000000000100100xx: _out=43;              //144-147
                32'b0000000000000000000000001001010x: _out=43;              //148-149
                
                32'b0000000000000000000000001001011x: _out=44;              //150-151
                32'b00000000000000000000000010011xxx: _out=44;              //152-159
                32'b00000000000000000000000010100xxx: _out=44;              //160-167
                
                32'b00000000000000000000000010101xxx: _out=45;              //168-175
                32'b00000000000000000000000010110xxx: _out=45;              //176-183
                32'b000000000000000000000000101110xx: _out=45;              //184-187
                32'b00000000000000000000000010111100: _out=45;              //188
                
                32'b00000000000000000000000010111101: _out=46;              //189
                32'b0000000000000000000000001011111x: _out=46;              //190-191
                32'b0000000000000000000000001100xxxx: _out=46;              //192-207
                32'b000000000000000000000000110100xx: _out=46;              //208-211
                
                32'b000000000000000000000000110101xx: _out=47;              //212-215
                32'b00000000000000000000000011011xxx: _out=47;              //216-223
                32'b00000000000000000000000011100xxx: _out=47;              //224-231
                32'b000000000000000000000000111010xx: _out=47;              //232-235
                32'b0000000000000000000000001110110x: _out=47;              //236-237
                
                32'b0000000000000000000000001110111x: _out=48;              //238-239
                32'b0000000000000000000000001111xxxx: _out=48;              //240-255
                32'b00000000000000000000000100000xxx: _out=48;              //256-263
                32'b0000000000000000000000010000100x: _out=48;              //264-265
                32'b00000000000000000000000100001010: _out=48;              //266
                
                32'b00000000000000000000000100001011: _out=49;              //267
                32'b000000000000000000000001000011xx: _out=49;              //268-271
                32'b0000000000000000000000010001xxxx: _out=49;              //272-287
                32'b00000000000000000000000100100xxx: _out=49;              //288-295
                32'b0000000000000000000000010010100x: _out=49;              //296-297
                32'b00000000000000000000000100101010: _out=49;              //298
                
                32'b00000000000000000000000100101011: _out=50;              //299
                32'b000000000000000000000001001011xx: _out=50;              //300-303
                32'b0000000000000000000000010011xxxx: _out=50;              //304-319
                32'b00000000000000000000000101000xxx: _out=50;              //320-327
                32'b000000000000000000000001010010xx: _out=50;              //328-331
                32'b0000000000000000000000010100110x: _out=50;              //332-333
                32'b00000000000000000000000101001110: _out=50;              //334
                
                32'b00000000000000000000000101001111: _out=51;              //335
                32'b0000000000000000000000010101xxxx: _out=51;              //336-351
                32'b0000000000000000000000010110xxxx: _out=51;              //352-367
                32'b00000000000000000000000101110xxx: _out=51;              //368-375
                
                32'b00000000000000000000000101111xxx: _out=52;              //376-383
                32'b000000000000000000000001100xxxxx: _out=52;              //384-415
                32'b000000000000000000000001101000xx: _out=52;              //416-419
                32'b0000000000000000000000011010010x: _out=52;              //420-421
                
                32'b0000000000000000000000011010011x: _out=53;              //422-423
                32'b00000000000000000000000110101xxx: _out=53;              //424-431
                32'b0000000000000000000000011011xxxx: _out=53;              //432-447
                32'b0000000000000000000000011100xxxx: _out=53;              //448-463
                32'b00000000000000000000000111010xxx: _out=53;              //464-471
                32'b0000000000000000000000011101100x: _out=53;              //472-473
                
                32'b0000000000000000000000011101101x: _out=54;              //474-475
                32'b000000000000000000000001110111xx: _out=54;              //476-479
                32'b000000000000000000000001111xxxxx: _out=54;              //480-511
                32'b0000000000000000000000100000xxxx: _out=54;              //512-527
                32'b0000000000000000000000100001000x: _out=54;              //528-529
                32'b00000000000000000000001000010010: _out=54;              //530
                
                32'b00000000000000000000001000010011: _out=55;              //531
                32'b000000000000000000000010000101xx: _out=55;              //532-535
                32'b00000000000000000000001000011xxx: _out=55;              //536-543
                32'b000000000000000000000010001xxxxx: _out=55;              //544-575
                32'b0000000000000000000000100100xxxx: _out=55;              //576-591
                32'b000000000000000000000010010100xx: _out=55;              //592-595
                
                32'b000000000000000000000010010101xx: _out=56;              //596-599
                32'b00000000000000000000001001011xxx: _out=56;              //600-607
                32'b000000000000000000000010011xxxxx: _out=56;              //608-639
                32'b0000000000000000000000101000xxxx: _out=56;              //640-655
                32'b00000000000000000000001010010xxx: _out=56;              //656-663
                32'b000000000000000000000010100110xx: _out=56;              //664-667
                32'b00000000000000000000001010011100: _out=56;              //668
                
                32'b00000000000000000000001010011101: _out=57;              //669
                32'b0000000000000000000000101001111x: _out=57;              //670-671
                32'b000000000000000000000010101xxxxx: _out=57;              //672-703
                32'b000000000000000000000010110xxxxx: _out=57;              //704-735
                32'b00000000000000000000001011100xxx: _out=57;              //736-743
                32'b000000000000000000000010111010xx: _out=57;              //744-747
                32'b0000000000000000000000101110110x: _out=57;              //748-749
                
                32'b0000000000000000000000101110111x: _out=58;              //750-751
                32'b0000000000000000000000101111xxxx: _out=58;              //752-767
                32'b00000000000000000000001100xxxxxx: _out=58;              //768-831
                32'b00000000000000000000001101000xxx: _out=58;              //832-839
                32'b0000000000000000000000110100100x: _out=58;              //840-841
                
                32'b0000000000000000000000110100101x: _out=59;              //842-843
                32'b000000000000000000000011010011xx: _out=59;              //844-847
                32'b0000000000000000000000110101xxxx: _out=59;              //848-863
                32'b000000000000000000000011011xxxxx: _out=59;              //864-895
                32'b000000000000000000000011100xxxxx: _out=59;              //896-927
                32'b0000000000000000000000111010xxxx: _out=59;              //928-943
                32'b00000000000000000000001110110000: _out=59;              //944
                
                32'b00000000000000000000001110110001: _out=60;              //945
                32'b0000000000000000000000111011001x: _out=60;              //946-947
                32'b000000000000000000000011101101xx: _out=60;              //948-951
                32'b00000000000000000000001110111xxx: _out=60;              //952-959
                32'b00000000000000000000001111xxxxxx: _out=60;              //960-1023
                32'b000000000000000000000100000xxxxx: _out=60;              //1024-1055
                32'b000000000000000000000100001000xx: _out=60;              //1056-1059
                
                32'b000000000000000000000100001001xx: _out=61;              //1060-1063
                32'b00000000000000000000010000101xxx: _out=61;              //1064-1071
                32'b0000000000000000000001000011xxxx: _out=61;              //1072-1087
                32'b00000000000000000000010001xxxxxx: _out=61;              //1088-1151
                32'b000000000000000000000100100xxxxx: _out=61;              //1152-1183
                32'b000000000000000000000100101000xx: _out=61;              //1184-1187
                32'b00000000000000000000010010100100: _out=61;              //1188
                
                32'b00000000000000000000010010100101: _out=62;              //1189
                32'b0000000000000000000001001010011x: _out=62;              //1190-1191
                32'b00000000000000000000010010101xxx: _out=62;              //1192-1199
                32'b0000000000000000000001001011xxxx: _out=62;              //1200-1215
                32'b00000000000000000000010011xxxxxx: _out=62;              //1216-1279
                32'b000000000000000000000101000xxxxx: _out=62;              //1280-1311
                32'b0000000000000000000001010010xxxx: _out=62;              //1312-1327
                32'b000000000000000000000101001100xx: _out=62;              //1328-1331
                32'b0000000000000000000001010011010x: _out=62;              //1332-1333
                
                32'b0000000000000000000001010011011x: _out=63;              //1334-1335
                32'b00000000000000000000010100111xxx: _out=63;              //1336-1343
                32'b00000000000000000000010101xxxxxx: _out=63;              //1344-1407
                32'b00000000000000000000010110xxxxxx: _out=63;              //1408-1471
                32'b0000000000000000000001011100xxxx: _out=63;              //1472-1487
                32'b00000000000000000000010111010xxx: _out=63;              //1488-1495
                32'b00000000000000000000010111011000: _out=63;              //1496
                
                32'b00000000000000000000010111011001: _out=64;              //1497
                32'b0000000000000000000001011101101x: _out=64;              //1498-1499
                32'b000000000000000000000101110111xx: _out=64;              //1500-1503
                32'b000000000000000000000101111xxxxx: _out=64;              //1504-1535
                32'b0000000000000000000001100xxxxxxx: _out=64;              //1536-1663
                32'b00000000000000000000011010000xxx: _out=64;              //1664-1671
                32'b000000000000000000000110100010xx: _out=64;              //1672-1675
                32'b0000000000000000000001101000110x: _out=64;              //1676-1677
                32'b00000000000000000000011010001110: _out=64;              //1678
                
                32'b00000000000000000000011010001111: _out=65;              //1679
                32'b0000000000000000000001101001xxxx: _out=65;              //1680-1695
                32'b000000000000000000000110101xxxxx: _out=65;              //1696-1727
                32'b00000000000000000000011011xxxxxx: _out=65;              //1728-1791
                32'b00000000000000000000011100xxxxxx: _out=65;              //1792-1855
                32'b0000000000000000000001110100xxxx: _out=65;              //1856-1871
                32'b00000000000000000000011101010xxx: _out=65;              //1872-1879
                32'b000000000000000000000111010110xx: _out=65;              //1880-1883
                
                32'b000000000000000000000111010111xx: _out=66;              //1884-1887
                32'b000000000000000000000111011xxxxx: _out=66;              //1888-1919
                32'b0000000000000000000001111xxxxxxx: _out=66;              //1920-2047
                32'b00000000000000000000100000xxxxxx: _out=66;              //2048-2111
                32'b0000000000000000000010000100000x: _out=66;              //2112-2113
                
                32'b0000000000000000000010000100001x: _out=67;              //2114-2115
                32'b000000000000000000001000010001xx: _out=67;              //2116-2119
                32'b00000000000000000000100001001xxx: _out=67;              //2120-2127
                32'b0000000000000000000010000101xxxx: _out=67;              //2128-2143
                32'b000000000000000000001000011xxxxx: _out=67;              //2144-2175
                32'b0000000000000000000010001xxxxxxx: _out=67;              //2176-2303
                32'b00000000000000000000100100xxxxxx: _out=67;              //2304-2367
                32'b000000000000000000001001010000xx: _out=67;              //2368-2371
                
                32'b000000000000000000001001010001xx: _out=68;              //2372-2375
                32'b00000000000000000000100101001xxx: _out=68;              //2376-2383
                32'b0000000000000000000010010101xxxx: _out=68;              //2384-2399
                32'b000000000000000000001001011xxxxx: _out=68;              //2400-2431
                32'b0000000000000000000010011xxxxxxx: _out=68;              //2432-2559
                32'b00000000000000000000101000xxxxxx: _out=68;              //2560-2623
                32'b000000000000000000001010010xxxxx: _out=68;              //2624-2655
                32'b000000000000000000001010011000xx: _out=68;              //2656-2659
                32'b00000000000000000000101001100100: _out=68;              //2660
                
                32'b00000000000000000000101001100101: _out=69;              //2661
                32'b0000000000000000000010100110011x: _out=69;              //2662-2663
                32'b00000000000000000000101001101xxx: _out=69;              //2664-2671
                32'b0000000000000000000010100111xxxx: _out=69;              //2672-2687
                32'b0000000000000000000010101xxxxxxx: _out=69;              //2688-2815
                32'b0000000000000000000010110xxxxxxx: _out=69;              //2816-2943
                32'b000000000000000000001011100xxxxx: _out=69;              //2944-2975
                32'b00000000000000000000101110100xxx: _out=69;              //2976-2983
                32'b0000000000000000000010111010100x: _out=69;              //2984-2985
                
                32'b0000000000000000000010111010101x: _out=70;              //2986-2987
                32'b000000000000000000001011101011xx: _out=70;              //2988-2991
                32'b0000000000000000000010111011xxxx: _out=70;              //2992-3007
                32'b00000000000000000000101111xxxxxx: _out=70;              //3008-3071
                32'b000000000000000000001100xxxxxxxx: _out=70;              //3072-3327
                32'b0000000000000000000011010000xxxx: _out=70;              //3328-3343
                32'b000000000000000000001101000100xx: _out=70;              //3344-3347
                32'b0000000000000000000011010001010x: _out=70;              //3348-3349
                
                32'b0000000000000000000011010001011x: _out=71;              //3350-3351
                32'b00000000000000000000110100011xxx: _out=71;              //3352-3359
                32'b000000000000000000001101001xxxxx: _out=71;              //3360-3391
                32'b00000000000000000000110101xxxxxx: _out=71;              //3392-3455
                32'b0000000000000000000011011xxxxxxx: _out=71;              //3456-3583
                32'b0000000000000000000011100xxxxxxx: _out=71;              //3584-3711
                32'b000000000000000000001110100xxxxx: _out=71;              //3712-3743
                32'b00000000000000000000111010100xxx: _out=71;              //3744-3751
                32'b000000000000000000001110101010xx: _out=71;              //3752-3755
                32'b0000000000000000000011101010110x: _out=71;              //3756-3757
                32'b00000000000000000000111010101110: _out=71;              //3758
                
                32'b00000000000000000000111010101111: _out=72;              //3759
                32'b0000000000000000000011101011xxxx: _out=72;              //3760-3775
                32'b00000000000000000000111011xxxxxx: _out=72;              //3776-3839
                32'b000000000000000000001111xxxxxxxx: _out=72;              //3840-4095
                32'b00000000000000000001000000xxxxxx: _out=72;              //4096-4159
                32'b000000000000000000010000010xxxxx: _out=72;              //4160-4191
                32'b0000000000000000000100000110xxxx: _out=72;              //4192-4207
                32'b00000000000000000001000001110xxx: _out=72;              //4208-4215
                32'b00000000000000000001000001111000: _out=72;              //4216
                
                32'b00000000000000000001000001111001: _out=73;              //4217
                32'b0000000000000000000100000111101x: _out=73;              //4218-4219
                32'b000000000000000000010000011111xx: _out=73;              //4220-4223
                32'b0000000000000000000100001xxxxxxx: _out=73;              //4224-4351
                32'b000000000000000000010001xxxxxxxx: _out=73;              //4352-4607
                32'b00000000000000000001001000xxxxxx: _out=73;              //4608-4671
                32'b000000000000000000010010010xxxxx: _out=73;              //4672-4703
                32'b0000000000000000000100100110xxxx: _out=73;              //4704-4719
                32'b00000000000000000001001001110xxx: _out=73;              //4720-4727
                32'b000000000000000000010010011110xx: _out=73;              //4728-4731
                
                32'b000000000000000000010010011111xx: _out=74;              //4732-4735
                32'b0000000000000000000100101xxxxxxx: _out=74;              //4736-4863
                32'b000000000000000000010011xxxxxxxx: _out=74;              //4864-5119
                32'b0000000000000000000101000xxxxxxx: _out=74;              //5120-5247
                32'b000000000000000000010100100xxxxx: _out=74;              //5248-5279
                32'b0000000000000000000101001010xxxx: _out=74;              //5280-5295
                32'b00000000000000000001010010110xxx: _out=74;              //5296-5303
                32'b000000000000000000010100101110xx: _out=74;              //5304-5307
                32'b00000000000000000001010010111100: _out=74;              //5308
                
                32'b00000000000000000001010010111101: _out=75;              //5309
                32'b0000000000000000000101001011111x: _out=75;              //5310-5311
                32'b00000000000000000001010011xxxxxx: _out=75;              //5312-5375
                32'b000000000000000000010101xxxxxxxx: _out=75;              //5376-5631
                32'b000000000000000000010110xxxxxxxx: _out=75;              //5632-5887
                32'b00000000000000000001011100xxxxxx: _out=75;              //5888-5951
                32'b000000000000000000010111010000xx: _out=75;              //5952-5955
                32'b00000000000000000001011101000100: _out=75;              //5956
                
                32'b00000000000000000001011101000101: _out=76;              //5957
                32'b0000000000000000000101110100011x: _out=76;              //5958-5959
                32'b00000000000000000001011101001xxx: _out=76;              //5960-5967
                32'b0000000000000000000101110101xxxx: _out=76;              //5968-5983
                32'b000000000000000000010111011xxxxx: _out=76;              //5984-6015
                32'b0000000000000000000101111xxxxxxx: _out=76;              //6016-6143
                32'b00000000000000000001100xxxxxxxxx: _out=76;              //6144-6655
                32'b0000000000000000000110100000xxxx: _out=76;              //6656-6671
                32'b00000000000000000001101000010xxx: _out=76;              //6672-6679
                32'b000000000000000000011010000110xx: _out=76;              //6680-6683
                
                32'b000000000000000000011010000111xx: _out=77;              //6684-6687
                32'b000000000000000000011010001xxxxx: _out=77;              //6688-6719
                32'b00000000000000000001101001xxxxxx: _out=77;              //6720-6783
                32'b0000000000000000000110101xxxxxxx: _out=77;              //6784-6911
                32'b000000000000000000011011xxxxxxxx: _out=77;              //6912-7167
                32'b000000000000000000011100xxxxxxxx: _out=77;              //7168-7423
                32'b00000000000000000001110100xxxxxx: _out=77;              //7424-7487
                32'b00000000000000000001110101000xxx: _out=77;              //7488-7495
                32'b0000000000000000000111010100100x: _out=77;              //7496-7497
                32'b00000000000000000001110101001010: _out=77;              //7498
                
                32'b00000000000000000001110101001011: _out=78;              //7499
                32'b000000000000000000011101010011xx: _out=78;              //7500-7503
                32'b0000000000000000000111010101xxxx: _out=78;              //7504-7519
                32'b000000000000000000011101011xxxxx: _out=78;              //7520-7551
                32'b0000000000000000000111011xxxxxxx: _out=78;              //7552-7679
                32'b00000000000000000001111xxxxxxxxx: _out=78;              //7680-8191
                32'b0000000000000000001000000xxxxxxx: _out=78;              //8192-8319
                32'b00000000000000000010000010xxxxxx: _out=78;              //8320-8383
                32'b0000000000000000001000001100xxxx: _out=78;              //8384-8399
                32'b00000000000000000010000011010xxx: _out=78;              //8400-8407
                32'b000000000000000000100000110110xx: _out=78;              //8408-8411
                32'b0000000000000000001000001101110x: _out=78;              //8412-8413
                
                32'b0000000000000000001000001101111x: _out=79;              //8414-8415
                32'b000000000000000000100000111xxxxx: _out=79;              //8416-8447
                32'b000000000000000000100001xxxxxxxx: _out=79;              //8448-8703
                32'b00000000000000000010001xxxxxxxxx: _out=79;              //8704-9215
                32'b0000000000000000001001000xxxxxxx: _out=79;              //9216-9343
                32'b00000000000000000010010010xxxxxx: _out=79;              //9344-9407
                32'b000000000000000000100100110xxxxx: _out=79;              //9408-9439
                32'b00000000000000000010010011100000: _out=79;              //9440
                
                32'b00000000000000000010010011100001: _out=80;              //9441
                32'b0000000000000000001001001110001x: _out=80;              //9442-9443
                32'b000000000000000000100100111001xx: _out=80;              //9444-9447
                32'b00000000000000000010010011101xxx: _out=80;              //9448-9455
                32'b0000000000000000001001001111xxxx: _out=80;              //9456-9471
                32'b000000000000000000100101xxxxxxxx: _out=80;              //9472-9727
                32'b00000000000000000010011xxxxxxxxx: _out=80;              //9728-10239
                32'b000000000000000000101000xxxxxxxx: _out=80;              //10240-10495
                32'b00000000000000000010100100xxxxxx: _out=80;              //10496-10559
                32'b000000000000000000101001010xxxxx: _out=80;              //10560-10591
                32'b00000000000000000010100101100000: _out=80;              //10592
                
                32'b00000000000000000010100101100001: _out=81;              //10593
                32'b0000000000000000001010010110001x: _out=81;              //10594-10595
                32'b000000000000000000101001011001xx: _out=81;              //10596-10599
                32'b00000000000000000010100101101xxx: _out=81;              //10600-10607
                32'b0000000000000000001010010111xxxx: _out=81;              //10608-10623
                32'b0000000000000000001010011xxxxxxx: _out=81;              //10624-10751
                32'b00000000000000000010101xxxxxxxxx: _out=81;              //10752-11263
                32'b00000000000000000010110xxxxxxxxx: _out=81;              //11264-11775
                32'b00000000000000000010111000xxxxxx: _out=81;              //11776-11839
                32'b000000000000000000101110010xxxxx: _out=81;              //11840-11871
                32'b00000000000000000010111001100xxx: _out=81;              //11872-11879
                32'b000000000000000000101110011010xx: _out=81;              //11880-11883
                32'b0000000000000000001011100110110x: _out=81;              //11884-11885
                
                32'b0000000000000000001011100110111x: _out=82;              //11886-11887
                32'b0000000000000000001011100111xxxx: _out=82;              //11888-11903
                32'b0000000000000000001011101xxxxxxx: _out=82;              //11904-12031
                32'b000000000000000000101111xxxxxxxx: _out=82;              //12032-12287
                32'b0000000000000000001100xxxxxxxxxx: _out=82;              //12288-13311
                32'b0000000000000000001101000000xxxx: _out=82;              //13312-13327
                32'b00000000000000000011010000010xxx: _out=82;              //13328-13335
                
                32'b00000000000000000011010000011xxx: _out=83;              //13336-13343
                32'b000000000000000000110100001xxxxx: _out=83;              //13344-13375
                32'b00000000000000000011010001xxxxxx: _out=83;              //13376-13439
                32'b0000000000000000001101001xxxxxxx: _out=83;              //13440-13567
                32'b000000000000000000110101xxxxxxxx: _out=83;              //13568-13823
                32'b00000000000000000011011xxxxxxxxx: _out=83;              //13824-14335
                32'b00000000000000000011100xxxxxxxxx: _out=83;              //14336-14847
                32'b00000000000000000011101000xxxxxx: _out=83;              //14848-14911
                32'b000000000000000000111010010xxxxx: _out=83;              //14912-14943
                32'b0000000000000000001110100110xxxx: _out=83;              //14944-14959
                32'b0000000000000000001110100111000x: _out=83;              //14960-14961
                32'b00000000000000000011101001110010: _out=83;              //14962
                
                32'b00000000000000000011101001110011: _out=84;              //14963
                32'b000000000000000000111010011101xx: _out=84;              //14964-14967
                32'b00000000000000000011101001111xxx: _out=84;              //14968-14975
                32'b0000000000000000001110101xxxxxxx: _out=84;              //14976-15103
                32'b000000000000000000111011xxxxxxxx: _out=84;              //15104-15359
                32'b0000000000000000001111xxxxxxxxxx: _out=84;              //15360-16383
                32'b000000000000000001000000xxxxxxxx: _out=84;              //16384-16639
                32'b0000000000000000010000010xxxxxxx: _out=84;              //16640-16767
                32'b0000000000000000010000011000xxxx: _out=84;              //16768-16783
                32'b000000000000000001000001100100xx: _out=84;              //16784-16787
                32'b00000000000000000100000110010100: _out=84;              //16788
                
                32'b00000000000000000100000110010101: _out=85;              //16789
                32'b0000000000000000010000011001011x: _out=85;              //16790-16791
                32'b00000000000000000100000110011xxx: _out=85;              //16792-16799
                32'b000000000000000001000001101xxxxx: _out=85;              //16800-16831
                32'b00000000000000000100000111xxxxxx: _out=85;              //16832-16895
                32'b00000000000000000100001xxxxxxxxx: _out=85;              //16896-17407
                32'b0000000000000000010001xxxxxxxxxx: _out=85;              //17408-18431
                32'b000000000000000001001000xxxxxxxx: _out=85;              //18432-18687
                32'b0000000000000000010010010xxxxxxx: _out=85;              //18688-18815
                32'b0000000000000000010010011000xxxx: _out=85;              //18816-18831
                32'b000000000000000001001001100100xx: _out=85;              //18832-18835
                32'b00000000000000000100100110010100: _out=85;              //18836
                
                32'b00000000000000000100100110010101: _out=86;              //18837
                32'b0000000000000000010010011001011x: _out=86;              //18838-18839
                32'b00000000000000000100100110011xxx: _out=86;              //18840-18847
                32'b000000000000000001001001101xxxxx: _out=86;              //18848-18879
                32'b00000000000000000100100111xxxxxx: _out=86;              //18880-18943
                32'b00000000000000000100101xxxxxxxxx: _out=86;              //18944-19455
                32'b0000000000000000010011xxxxxxxxxx: _out=86;              //19456-20479
                32'b00000000000000000101000xxxxxxxxx: _out=86;              //20480-20991
                32'b0000000000000000010100100xxxxxxx: _out=86;              //20992-21119
                32'b00000000000000000101001010000xxx: _out=86;              //21120-21127
                32'b000000000000000001010010100010xx: _out=86;              //21128-21131
                32'b0000000000000000010100101000110x: _out=86;              //21132-21133
                32'b00000000000000000101001010001110: _out=86;              //21134
                
                32'b00000000000000000101001010001111: _out=87;              //21135
                32'b0000000000000000010100101001xxxx: _out=87;              //21136-21151
                32'b000000000000000001010010101xxxxx: _out=87;              //21152-21183
                32'b00000000000000000101001011xxxxxx: _out=87;              //21184-21247
                32'b000000000000000001010011xxxxxxxx: _out=87;              //21248-21503
                32'b0000000000000000010101xxxxxxxxxx: _out=87;              //21504-22527
                32'b0000000000000000010110xxxxxxxxxx: _out=87;              //22528-23551
                32'b0000000000000000010111000xxxxxxx: _out=87;              //23552-23679
                32'b000000000000000001011100100xxxxx: _out=87;              //23680-23711
                32'b0000000000000000010111001010000x: _out=87;              //23712-23713
                
                32'b0000000000000000010111001010001x: _out=88;              //23714-23715
                32'b000000000000000001011100101001xx: _out=88;              //23716-23719
                32'b00000000000000000101110010101xxx: _out=88;              //23720-23727
                32'b0000000000000000010111001011xxxx: _out=88;              //23728-23743
                32'b00000000000000000101110011xxxxxx: _out=88;              //23744-23807
                32'b000000000000000001011101xxxxxxxx: _out=88;              //23808-24063
                32'b00000000000000000101111xxxxxxxxx: _out=88;              //24064-24575
                32'b0000000000000000011000xxxxxxxxxx: _out=88;              //24576-25599
                32'b00000000000000000110010xxxxxxxxx: _out=88;              //25600-26111
                32'b000000000000000001100110xxxxxxxx: _out=88;              //26112-26367
                32'b0000000000000000011001110xxxxxxx: _out=88;              //26368-26495
                32'b00000000000000000110011110xxxxxx: _out=88;              //26496-26559
                32'b000000000000000001100111110xxxxx: _out=88;              //26560-26591
                32'b0000000000000000011001111110xxxx: _out=88;              //26592-26607
                
                32'b0000000000000000011001111111xxxx: _out=89;              //26608-26623
                32'b000000000000000001101xxxxxxxxxxx: _out=89;              //26624-28671
                32'b0000000000000000011100xxxxxxxxxx: _out=89;              //28672-29695
                32'b0000000000000000011101000xxxxxxx: _out=89;              //29696-29823
                32'b0000000000000000011101001000xxxx: _out=89;              //29824-29839
                32'b00000000000000000111010010010xxx: _out=89;              //29840-29847
                32'b000000000000000001110100100110xx: _out=89;              //29848-29851
                32'b0000000000000000011101001001110x: _out=89;              //29852-29853
                
                32'b0000000000000000011101001001111x: _out=90;              //29854-29855
                32'b000000000000000001110100101xxxxx: _out=90;              //29856-29887
                32'b00000000000000000111010011xxxxxx: _out=90;              //29888-29951
                32'b000000000000000001110101xxxxxxxx: _out=90;              //29952-30207
                32'b00000000000000000111011xxxxxxxxx: _out=90;              //30208-30719
                32'b000000000000000001111xxxxxxxxxxx: _out=90;              //30720-32767
                32'b00000000000000001000000xxxxxxxxx: _out=90;              //32768-33279
                32'b0000000000000000100000100xxxxxxx: _out=90;              //33280-33407
                32'b00000000000000001000001010xxxxxx: _out=90;              //33408-33471
                32'b0000000000000000100000101100xxxx: _out=90;              //33472-33487
                32'b00000000000000001000001011010xxx: _out=90;              //33488-33495
                32'b00000000000000001000001011011000: _out=90;              //33496
                
                32'b00000000000000001000001011011001: _out=91;              //33497
                32'b0000000000000000100000101101101x: _out=91;              //33498-33499
                32'b000000000000000010000010110111xx: _out=91;              //33500-33503
                32'b000000000000000010000010111xxxxx: _out=91;              //33504-33535
                32'b000000000000000010000011xxxxxxxx: _out=91;              //33536-33791
                32'b0000000000000000100001xxxxxxxxxx: _out=91;              //33792-34815
                32'b000000000000000010001xxxxxxxxxxx: _out=91;              //34816-36863
                32'b00000000000000001001000xxxxxxxxx: _out=91;              //36864-37375
                32'b0000000000000000100100100xxxxxxx: _out=91;              //37376-37503
                32'b00000000000000001001001010xxxxxx: _out=91;              //37504-37567
                32'b0000000000000000100100101100xxxx: _out=91;              //37568-37583
                
                32'b0000000000000000100100101101xxxx: _out=92;              //37584-37599
                32'b000000000000000010010010111xxxxx: _out=92;              //37600-37631
                32'b000000000000000010010011xxxxxxxx: _out=92;              //37632-37887
                32'b0000000000000000100101xxxxxxxxxx: _out=92;              //37888-38911
                32'b000000000000000010011xxxxxxxxxxx: _out=92;              //38912-40959
                32'b0000000000000000101000xxxxxxxxxx: _out=92;              //40960-41983
                32'b0000000000000000101001000xxxxxxx: _out=92;              //41984-42111
                32'b000000000000000010100100100xxxxx: _out=92;              //42112-42143
                32'b0000000000000000101001001010xxxx: _out=92;              //42144-42159
                32'b00000000000000001010010010110xxx: _out=92;              //42160-42167
                32'b0000000000000000101001001011100x: _out=92;              //42168-42169
                
                32'b0000000000000000101001001011101x: _out=93;              //42170-42171
                32'b000000000000000010100100101111xx: _out=93;              //42172-42175
                32'b00000000000000001010010011xxxxxx: _out=93;              //42176-42239
                32'b000000000000000010100101xxxxxxxx: _out=93;              //42240-42495
                32'b00000000000000001010011xxxxxxxxx: _out=93;              //42496-43007
                32'b000000000000000010101xxxxxxxxxxx: _out=93;              //43008-45055
                32'b000000000000000010110xxxxxxxxxxx: _out=93;              //45056-47103
                32'b0000000000000000101110000xxxxxxx: _out=93;              //47104-47231
                32'b00000000000000001011100010xxxxxx: _out=93;              //47232-47295
                32'b0000000000000000101110001100xxxx: _out=93;              //47296-47311
                32'b000000000000000010111000110100xx: _out=93;              //47312-47315
                
                32'b000000000000000010111000110101xx: _out=94;              //47316-47319
                32'b00000000000000001011100011011xxx: _out=94;              //47320-47327
                32'b000000000000000010111000111xxxxx: _out=94;              //47328-47359
                32'b000000000000000010111001xxxxxxxx: _out=94;              //47360-47615
                32'b00000000000000001011101xxxxxxxxx: _out=94;              //47616-48127
                32'b0000000000000000101111xxxxxxxxxx: _out=94;              //48128-49151
                32'b000000000000000011000xxxxxxxxxxx: _out=94;              //49152-51199
                32'b0000000000000000110010xxxxxxxxxx: _out=94;              //51200-52223
                32'b00000000000000001100110xxxxxxxxx: _out=94;              //52224-52735
                32'b000000000000000011001110xxxxxxxx: _out=94;              //52736-52991
                32'b00000000000000001100111100xxxxxx: _out=94;              //52992-53055
                32'b000000000000000011001111010xxxxx: _out=94;              //53056-53087
                32'b00000000000000001100111101100000: _out=94;              //53088
                
                32'b00000000000000001100111101100001: _out=95;              //53089
                32'b0000000000000000110011110110001x: _out=95;              //53090-53091
                32'b000000000000000011001111011001xx: _out=95;              //53092-53095
                32'b00000000000000001100111101101xxx: _out=95;              //53096-53103
                32'b0000000000000000110011110111xxxx: _out=95;              //53104-53119
                32'b0000000000000000110011111xxxxxxx: _out=95;              //53120-53247
                32'b00000000000000001101xxxxxxxxxxxx: _out=95;              //53248-57343
                32'b000000000000000011100xxxxxxxxxxx: _out=95;              //57344-59391
                32'b0000000000000000111010000xxxxxxx: _out=95;              //59392-59519
                32'b000000000000000011101000100xxxxx: _out=95;              //59520-59551
                32'b00000000000000001110100010100xxx: _out=95;              //59552-59559
                32'b000000000000000011101000101010xx: _out=95;              //59560-59563
                32'b0000000000000000111010001010110x: _out=95;              //59564-59565
                32'b00000000000000001110100010101110: _out=95;              //59566
                
                32'b00000000000000001110100010101111: _out=96;              //59567
                32'b0000000000000000111010001011xxxx: _out=96;              //59568-59583
                32'b00000000000000001110100011xxxxxx: _out=96;              //59584-59647
                32'b000000000000000011101001xxxxxxxx: _out=96;              //59648-59903
                32'b00000000000000001110101xxxxxxxxx: _out=96;              //59904-60415
                32'b0000000000000000111011xxxxxxxxxx: _out=96;              //60416-61439
                32'b00000000000000001111xxxxxxxxxxxx: _out=96;              //61440-65535
                32'b0000000000000001000000xxxxxxxxxx: _out=96;              //65536-66559
                32'b000000000000000100000100xxxxxxxx: _out=96;              //66560-66815
                32'b0000000000000001000001010000xxxx: _out=96;              //66816-66831
                32'b0000000000000001000001010001000x: _out=96;              //66832-66833
                32'b00000000000000010000010100010010: _out=96;              //66834
                
                32'b00000000000000010000010100010011: _out=97;              //66835
                32'b000000000000000100000101000101xx: _out=97;              //66836-66839
                32'b00000000000000010000010100011xxx: _out=97;              //66840-66847
                32'b000000000000000100000101001xxxxx: _out=97;              //66848-66879
                32'b00000000000000010000010101xxxxxx: _out=97;              //66880-66943
                32'b0000000000000001000001011xxxxxxx: _out=97;              //66944-67071
                32'b00000000000000010000011xxxxxxxxx: _out=97;              //67072-67583
                32'b000000000000000100001xxxxxxxxxxx: _out=97;              //67584-69631
                32'b00000000000000010001xxxxxxxxxxxx: _out=97;              //69632-73727
                32'b0000000000000001001000xxxxxxxxxx: _out=97;              //73728-74751
                32'b0000000000000001001001000xxxxxxx: _out=97;              //74752-74879
                32'b00000000000000010010010010xxxxxx: _out=97;              //74880-74943
                32'b000000000000000100100100110xxxxx: _out=97;              //74944-74975
                32'b00000000000000010010010011100xxx: _out=97;              //74976-74983
                32'b000000000000000100100100111010xx: _out=97;              //74984-74987
                32'b0000000000000001001001001110110x: _out=97;              //74988-74989
                
                32'b0000000000000001001001001110111x: _out=98;              //74990-74991
                32'b0000000000000001001001001111xxxx: _out=98;              //74992-75007
                32'b000000000000000100100101xxxxxxxx: _out=98;              //75008-75263
                32'b00000000000000010010011xxxxxxxxx: _out=98;              //75264-75775
                32'b000000000000000100101xxxxxxxxxxx: _out=98;              //75776-77823
                32'b00000000000000010011xxxxxxxxxxxx: _out=98;              //77824-81919
                32'b000000000000000101000xxxxxxxxxxx: _out=98;              //81920-83967
                32'b0000000000000001010010000xxxxxxx: _out=98;              //83968-84095
                32'b000000000000000101001000100xxxxx: _out=98;              //84096-84127
                32'b00000000000000010100100010100xxx: _out=98;              //84128-84135
                32'b000000000000000101001000101010xx: _out=98;              //84136-84139
                
                32'b000000000000000101001000101011xx: _out=99;              //84140-84143
                32'b0000000000000001010010001011xxxx: _out=99;              //84144-84159
                32'b00000000000000010100100011xxxxxx: _out=99;              //84160-84223
                32'b000000000000000101001001xxxxxxxx: _out=99;              //84224-84479
                32'b00000000000000010100101xxxxxxxxx: _out=99;              //84480-84991
                32'b0000000000000001010011xxxxxxxxxx: _out=99;              //84992-86015
                32'b00000000000000010101xxxxxxxxxxxx: _out=99;              //86016-90111
                32'b00000000000000010110xxxxxxxxxxxx: _out=99;              //90112-94207
                32'b0000000000000001011100000xxxxxxx: _out=99;              //94208-94335
                32'b00000000000000010111000010xxxxxx: _out=99;              //94336-94399
                32'b000000000000000101110000110000xx: _out=99;              //94400-94403
                32'b0000000000000001011100001100010x: _out=99;              //94404-94405
                32'b00000000000000010111000011000110: _out=99;              //94406
                
                32'b00000000000000010111000011000111: _out=100;              //94407
                32'b00000000000000010111000011001xxx: _out=100;              //94408-94415
                32'b0000000000000001011100001101xxxx: _out=100;              //94416-94431
                32'b000000000000000101110000111xxxxx: _out=100;              //94432-94463
                32'b000000000000000101110001xxxxxxxx: _out=100;              //94464-94719
                32'b00000000000000010111001xxxxxxxxx: _out=100;              //94720-95231
                32'b0000000000000001011101xxxxxxxxxx: _out=100;              //95232-96255
                32'b000000000000000101111xxxxxxxxxxx: _out=100;              //96256-98303
                32'b00000000000000011000xxxxxxxxxxxx: _out=100;              //98304-102399
                32'b000000000000000110010xxxxxxxxxxx: _out=100;              //102400-104447
                32'b0000000000000001100110xxxxxxxxxx: _out=100;              //104448-105471
                32'b000000000000000110011100xxxxxxxx: _out=100;              //105472-105727
                32'b0000000000000001100111010xxxxxxx: _out=100;              //105728-105855
                32'b00000000000000011001110110xxxxxx: _out=100;              //105856-105919
                32'b000000000000000110011101110000xx: _out=100;              //105920-105923
                32'b0000000000000001100111011100010x: _out=100;              //105924-105925
                
                32'b0000000000000001100111011100011x: _out=101;              //105926-105927
                32'b00000000000000011001110111001xxx: _out=101;              //105928-105935
                32'b0000000000000001100111011101xxxx: _out=101;              //105936-105951
                32'b000000000000000110011101111xxxxx: _out=101;              //105952-105983
                32'b00000000000000011001111xxxxxxxxx: _out=101;              //105984-106495
                32'b0000000000000001101xxxxxxxxxxxxx: _out=101;              //106496-114687
                32'b00000000000000011100xxxxxxxxxxxx: _out=101;              //114688-118783
                32'b00000000000000011101000000xxxxxx: _out=101;              //118784-118847
                32'b0000000000000001110100000100000x: _out=101;              //118848-118849
                32'b00000000000000011101000001000010: _out=101;              //118850
                
                32'b00000000000000011101000001000011: _out=102;              //118851
                32'b000000000000000111010000010001xx: _out=102;              //118852-118855
                32'b00000000000000011101000001001xxx: _out=102;              //118856-118863
                32'b0000000000000001110100000101xxxx: _out=102;              //118864-118879
                32'b000000000000000111010000011xxxxx: _out=102;              //118880-118911
                32'b0000000000000001110100001xxxxxxx: _out=102;              //118912-119039
                32'b000000000000000111010001xxxxxxxx: _out=102;              //119040-119295
                32'b00000000000000011101001xxxxxxxxx: _out=102;              //119296-119807
                32'b0000000000000001110101xxxxxxxxxx: _out=102;              //119808-120831
                32'b000000000000000111011xxxxxxxxxxx: _out=102;              //120832-122879
                32'b0000000000000001111xxxxxxxxxxxxx: _out=102;              //122880-131071
                32'b000000000000001000000xxxxxxxxxxx: _out=102;              //131072-133119
                32'b0000000000000010000010000xxxxxxx: _out=102;              //133120-133247
                32'b00000000000000100000100010xxxxxx: _out=102;              //133248-133311
                32'b000000000000001000001000110xxxxx: _out=102;              //133312-133343
                32'b00000000000000100000100011100xxx: _out=102;              //133344-133351
                32'b00000000000000100000100011101000: _out=102;              //133352
                
                32'b00000000000000100000100011101001: _out=103;              //133353
                32'b0000000000000010000010001110101x: _out=103;              //133354-133355
                32'b000000000000001000001000111011xx: _out=103;              //133356-133359
                32'b0000000000000010000010001111xxxx: _out=103;              //133360-133375
                32'b000000000000001000001001xxxxxxxx: _out=103;              //133376-133631
                32'b00000000000000100000101xxxxxxxxx: _out=103;              //133632-134143
                32'b0000000000000010000011xxxxxxxxxx: _out=103;              //134144-135167
                32'b00000000000000100001xxxxxxxxxxxx: _out=103;              //135168-139263
                32'b0000000000000010001xxxxxxxxxxxxx: _out=103;              //139264-147455
                32'b000000000000001001000xxxxxxxxxxx: _out=103;              //147456-149503
                32'b00000000000000100100100000xxxxxx: _out=103;              //149504-149567
                32'b000000000000001001001000010xxxxx: _out=103;              //149568-149599
                32'b0000000000000010010010000110xxxx: _out=103;              //149600-149615
                32'b00000000000000100100100001110xxx: _out=103;              //149616-149623
                
                32'b00000000000000100100100001111xxx: _out=104;              //149624-149631
                32'b0000000000000010010010001xxxxxxx: _out=104;              //149632-149759
                32'b000000000000001001001001xxxxxxxx: _out=104;              //149760-150015
                32'b00000000000000100100101xxxxxxxxx: _out=104;              //150016-150527
                32'b0000000000000010010011xxxxxxxxxx: _out=104;              //150528-151551
                32'b00000000000000100101xxxxxxxxxxxx: _out=104;              //151552-155647
                32'b0000000000000010011xxxxxxxxxxxxx: _out=104;              //155648-163839
                32'b000000000000001010000xxxxxxxxxxx: _out=104;              //163840-165887
                32'b0000000000000010100010xxxxxxxxxx: _out=104;              //165888-166911
                32'b00000000000000101000110xxxxxxxxx: _out=104;              //166912-167423
                32'b000000000000001010001110xxxxxxxx: _out=104;              //167424-167679
                32'b0000000000000010100011110xxxxxxx: _out=104;              //167680-167807
                32'b00000000000000101000111110xxxxxx: _out=104;              //167808-167871
                32'b00000000000000101000111111000xxx: _out=104;              //167872-167879
                32'b00000000000000101000111111001000: _out=104;              //167880
                
                32'b00000000000000101000111111001001: _out=105;              //167881
                32'b0000000000000010100011111100101x: _out=105;              //167882-167883
                32'b000000000000001010001111110011xx: _out=105;              //167884-167887
                32'b0000000000000010100011111101xxxx: _out=105;              //167888-167903
                32'b000000000000001010001111111xxxxx: _out=105;              //167904-167935
                32'b00000000000000101001xxxxxxxxxxxx: _out=105;              //167936-172031
                32'b0000000000000010101xxxxxxxxxxxxx: _out=105;              //172032-180223
                32'b00000000000000101100xxxxxxxxxxxx: _out=105;              //180224-184319
                32'b000000000000001011010xxxxxxxxxxx: _out=105;              //184320-186367
                32'b0000000000000010110110xxxxxxxxxx: _out=105;              //186368-187391
                32'b00000000000000101101110xxxxxxxxx: _out=105;              //187392-187903
                32'b000000000000001011011110xxxxxxxx: _out=105;              //187904-188159
                32'b0000000000000010110111110xxxxxxx: _out=105;              //188160-188287
                32'b00000000000000101101111110xxxxxx: _out=105;              //188288-188351
                32'b00000000000000101101111111000xxx: _out=105;              //188352-188359
                32'b000000000000001011011111110010xx: _out=105;              //188360-188363
                32'b00000000000000101101111111001100: _out=105;              //188364
                
                32'b00000000000000101101111111001101: _out=106;              //188365
                32'b0000000000000010110111111100111x: _out=106;              //188366-188367
                32'b0000000000000010110111111101xxxx: _out=106;              //188368-188383
                32'b000000000000001011011111111xxxxx: _out=106;              //188384-188415
                32'b0000000000000010111xxxxxxxxxxxxx: _out=106;              //188416-196607
                32'b0000000000000011000xxxxxxxxxxxxx: _out=106;              //196608-204799
                32'b00000000000000110010xxxxxxxxxxxx: _out=106;              //204800-208895
                32'b000000000000001100110xxxxxxxxxxx: _out=106;              //208896-210943
                32'b000000000000001100111000xxxxxxxx: _out=106;              //210944-211199
                32'b0000000000000011001110010xxxxxxx: _out=106;              //211200-211327
                32'b0000000000000011001110011000xxxx: _out=106;              //211328-211343
                32'b000000000000001100111001100100xx: _out=106;              //211344-211347
                32'b00000000000000110011100110010100: _out=106;              //211348
                
                32'b00000000000000110011100110010101: _out=107;              //211349
                32'b0000000000000011001110011001011x: _out=107;              //211350-211351
                32'b00000000000000110011100110011xxx: _out=107;              //211352-211359
                32'b000000000000001100111001101xxxxx: _out=107;              //211360-211391
                32'b00000000000000110011100111xxxxxx: _out=107;              //211392-211455
                32'b00000000000000110011101xxxxxxxxx: _out=107;              //211456-211967
                32'b0000000000000011001111xxxxxxxxxx: _out=107;              //211968-212991
                32'b000000000000001101xxxxxxxxxxxxxx: _out=107;              //212992-229375
                32'b00000000000000111000xxxxxxxxxxxx: _out=107;              //229376-233471
                32'b000000000000001110010xxxxxxxxxxx: _out=107;              //233472-235519
                32'b0000000000000011100110xxxxxxxxxx: _out=107;              //235520-236543
                32'b00000000000000111001110xxxxxxxxx: _out=107;              //236544-237055
                32'b00000000000000111001111000xxxxxx: _out=107;              //237056-237119
                32'b0000000000000011100111100100xxxx: _out=107;              //237120-237135
                32'b0000000000000011100111100101000x: _out=107;              //237136-237137
                
                32'b0000000000000011100111100101001x: _out=108;              //237138-237139
                32'b000000000000001110011110010101xx: _out=108;              //237140-237143
                32'b00000000000000111001111001011xxx: _out=108;              //237144-237151
                32'b000000000000001110011110011xxxxx: _out=108;              //237152-237183
                32'b0000000000000011100111101xxxxxxx: _out=108;              //237184-237311
                32'b000000000000001110011111xxxxxxxx: _out=108;              //237312-237567
                32'b0000000000000011101xxxxxxxxxxxxx: _out=108;              //237568-245759
                32'b000000000000001111xxxxxxxxxxxxxx: _out=108;              //245760-262143
                32'b000000000000010000000xxxxxxxxxxx: _out=108;              //262144-264191
                32'b0000000000000100000010xxxxxxxxxx: _out=108;              //264192-265215
                32'b00000000000001000000110xxxxxxxxx: _out=108;              //265216-265727
                32'b000000000000010000001110xxxxxxxx: _out=108;              //265728-265983
                32'b00000000000001000000111100xxxxxx: _out=108;              //265984-266047
                32'b0000000000000100000011110100xxxx: _out=108;              //266048-266063
                32'b00000000000001000000111101010xxx: _out=108;              //266064-266071
                32'b00000000000001000000111101011000: _out=108;              //266072
                
                32'b00000000000001000000111101011001: _out=109;              //266073
                32'b0000000000000100000011110101101x: _out=109;              //266074-266075
                32'b000000000000010000001111010111xx: _out=109;              //266076-266079
                32'b000000000000010000001111011xxxxx: _out=109;              //266080-266111
                32'b0000000000000100000011111xxxxxxx: _out=109;              //266112-266239
                32'b00000000000001000001xxxxxxxxxxxx: _out=109;              //266240-270335
                32'b0000000000000100001xxxxxxxxxxxxx: _out=109;              //270336-278527
                32'b000000000000010001xxxxxxxxxxxxxx: _out=109;              //278528-294911
                32'b000000000000010010000xxxxxxxxxxx: _out=109;              //294912-296959
                32'b0000000000000100100010xxxxxxxxxx: _out=109;              //296960-297983
                32'b00000000000001001000110xxxxxxxxx: _out=109;              //297984-298495
                32'b000000000000010010001110000xxxxx: _out=109;              //298496-298527
                32'b00000000000001001000111000100xxx: _out=109;              //298528-298535
                32'b0000000000000100100011100010100x: _out=109;              //298536-298537
                32'b00000000000001001000111000101010: _out=109;              //298538
                
                32'b00000000000001001000111000101011: _out=110;              //298539
                32'b000000000000010010001110001011xx: _out=110;              //298540-298543
                32'b0000000000000100100011100011xxxx: _out=110;              //298544-298559
                32'b00000000000001001000111001xxxxxx: _out=110;              //298560-298623
                32'b0000000000000100100011101xxxxxxx: _out=110;              //298624-298751
                32'b000000000000010010001111xxxxxxxx: _out=110;              //298752-299007
                32'b00000000000001001001xxxxxxxxxxxx: _out=110;              //299008-303103
                32'b0000000000000100101xxxxxxxxxxxxx: _out=110;              //303104-311295
                32'b000000000000010011xxxxxxxxxxxxxx: _out=110;              //311296-327679
                32'b00000000000001010000xxxxxxxxxxxx: _out=110;              //327680-331775
                32'b000000000000010100010xxxxxxxxxxx: _out=110;              //331776-333823
                32'b0000000000000101000110xxxxxxxxxx: _out=110;              //333824-334847
                32'b00000000000001010001110000xxxxxx: _out=110;              //334848-334911
                32'b000000000000010100011100010xxxxx: _out=110;              //334912-334943
                32'b0000000000000101000111000110xxxx: _out=110;              //334944-334959
                32'b000000000000010100011100011100xx: _out=110;              //334960-334963
                32'b0000000000000101000111000111010x: _out=110;              //334964-334965
                
                32'b0000000000000101000111000111011x: _out=111;              //334966-334967
                32'b00000000000001010001110001111xxx: _out=111;              //334968-334975
                32'b0000000000000101000111001xxxxxxx: _out=111;              //334976-335103
                32'b000000000000010100011101xxxxxxxx: _out=111;              //335104-335359
                32'b00000000000001010001111xxxxxxxxx: _out=111;              //335360-335871
                32'b0000000000000101001xxxxxxxxxxxxx: _out=111;              //335872-344063
                32'b000000000000010101xxxxxxxxxxxxxx: _out=111;              //344064-360447
                32'b0000000000000101100xxxxxxxxxxxxx: _out=111;              //360448-368639
                32'b00000000000001011010xxxxxxxxxxxx: _out=111;              //368640-372735
                32'b000000000000010110110xxxxxxxxxxx: _out=111;              //372736-374783
                32'b0000000000000101101110xxxxxxxxxx: _out=111;              //374784-375807
                32'b0000000000000101101111000000xxxx: _out=111;              //375808-375823
                32'b00000000000001011011110000010xxx: _out=111;              //375824-375831
                32'b000000000000010110111100000110xx: _out=111;              //375832-375835
                32'b0000000000000101101111000001110x: _out=111;              //375836-375837
                
                32'b0000000000000101101111000001111x: _out=112;              //375838-375839
                32'b000000000000010110111100001xxxxx: _out=112;              //375840-375871
                32'b00000000000001011011110001xxxxxx: _out=112;              //375872-375935
                32'b0000000000000101101111001xxxxxxx: _out=112;              //375936-376063
                32'b000000000000010110111101xxxxxxxx: _out=112;              //376064-376319
                32'b00000000000001011011111xxxxxxxxx: _out=112;              //376320-376831
                32'b000000000000010111xxxxxxxxxxxxxx: _out=112;              //376832-393215
                32'b000000000000011000xxxxxxxxxxxxxx: _out=112;              //393216-409599
                32'b0000000000000110010xxxxxxxxxxxxx: _out=112;              //409600-417791
                32'b000000000000011001100xxxxxxxxxxx: _out=112;              //417792-419839
                32'b0000000000000110011010xxxxxxxxxx: _out=112;              //419840-420863
                32'b00000000000001100110110xxxxxxxxx: _out=112;              //420864-421375
                32'b000000000000011001101110xxxxxxxx: _out=112;              //421376-421631
                32'b00000000000001100110111100xxxxxx: _out=112;              //421632-421695
                32'b00000000000001100110111101000000: _out=112;              //421696
                
                32'b00000000000001100110111101000001: _out=113;              //421697
                32'b0000000000000110011011110100001x: _out=113;              //421698-421699
                32'b000000000000011001101111010001xx: _out=113;              //421700-421703
                32'b00000000000001100110111101001xxx: _out=113;              //421704-421711
                32'b0000000000000110011011110101xxxx: _out=113;              //421712-421727
                32'b000000000000011001101111011xxxxx: _out=113;              //421728-421759
                32'b0000000000000110011011111xxxxxxx: _out=113;              //421760-421887
                32'b00000000000001100111xxxxxxxxxxxx: _out=113;              //421888-425983
                32'b00000000000001101xxxxxxxxxxxxxxx: _out=113;              //425984-458751
                32'b0000000000000111000xxxxxxxxxxxxx: _out=113;              //458752-466943
                32'b00000000000001110010xxxxxxxxxxxx: _out=113;              //466944-471039
                32'b000000000000011100110xxxxxxxxxxx: _out=113;              //471040-473087
                32'b00000000000001110011100000xxxxxx: _out=113;              //473088-473151
                
                32'b00000000000001110011100001xxxxxx: _out=114;              //473152-473215
                32'b0000000000000111001110001xxxxxxx: _out=114;              //473216-473343
                32'b000000000000011100111001xxxxxxxx: _out=114;              //473344-473599
                32'b00000000000001110011101xxxxxxxxx: _out=114;              //473600-474111
                32'b0000000000000111001111xxxxxxxxxx: _out=114;              //474112-475135
                32'b000000000000011101xxxxxxxxxxxxxx: _out=114;              //475136-491519
                32'b00000000000001111xxxxxxxxxxxxxxx: _out=114;              //491520-524287
                32'b00000000000010000000xxxxxxxxxxxx: _out=114;              //524288-528383
                32'b000000000000100000010xxxxxxxxxxx: _out=114;              //528384-530431
                32'b000000000000100000011000xxxxxxxx: _out=114;              //530432-530687
                32'b0000000000001000000110010xxxxxxx: _out=114;              //530688-530815
                32'b00000000000010000001100110xxxxxx: _out=114;              //530816-530879
                32'b000000000000100000011001110000xx: _out=114;              //530880-530883
                32'b00000000000010000001100111000100: _out=114;              //530884
                
                32'b00000000000010000001100111000101: _out=115;              //530885
                32'b0000000000001000000110011100011x: _out=115;              //530886-530887
                32'b00000000000010000001100111001xxx: _out=115;              //530888-530895
                32'b0000000000001000000110011101xxxx: _out=115;              //530896-530911
                32'b000000000000100000011001111xxxxx: _out=115;              //530912-530943
                32'b00000000000010000001101xxxxxxxxx: _out=115;              //530944-531455
                32'b0000000000001000000111xxxxxxxxxx: _out=115;              //531456-532479
                32'b0000000000001000001xxxxxxxxxxxxx: _out=115;              //532480-540671
                32'b000000000000100001xxxxxxxxxxxxxx: _out=115;              //540672-557055
                32'b00000000000010001xxxxxxxxxxxxxxx: _out=115;              //557056-589823
                32'b00000000000010010000xxxxxxxxxxxx: _out=115;              //589824-593919
                32'b0000000000001001000100xxxxxxxxxx: _out=115;              //593920-594943
                32'b00000000000010010001010xxxxxxxxx: _out=115;              //594944-595455
                32'b0000000000001001000101100xxxxxxx: _out=115;              //595456-595583
                32'b00000000000010010001011010xxxxxx: _out=115;              //595584-595647
                32'b00000000000010010001011011000xxx: _out=115;              //595648-595655
                32'b000000000000100100010110110010xx: _out=115;              //595656-595659
                32'b0000000000001001000101101100110x: _out=115;              //595660-595661
                32'b00000000000010010001011011001110: _out=115;              //595662
                
                32'b00000000000010010001011011001111: _out=116;              //595663
                32'b0000000000001001000101101101xxxx: _out=116;              //595664-595679
                32'b000000000000100100010110111xxxxx: _out=116;              //595680-595711
                32'b000000000000100100010111xxxxxxxx: _out=116;              //595712-595967
                32'b000000000000100100011xxxxxxxxxxx: _out=116;              //595968-598015
                32'b0000000000001001001xxxxxxxxxxxxx: _out=116;              //598016-606207
                32'b000000000000100101xxxxxxxxxxxxxx: _out=116;              //606208-622591
                32'b00000000000010011xxxxxxxxxxxxxxx: _out=116;              //622592-655359
                32'b0000000000001010000xxxxxxxxxxxxx: _out=116;              //655360-663551
                32'b00000000000010100010xxxxxxxxxxxx: _out=116;              //663552-667647
                32'b00000000000010100011000xxxxxxxxx: _out=116;              //667648-668159
                32'b0000000000001010001100100xxxxxxx: _out=116;              //668160-668287
                32'b000000000000101000110010100xxxxx: _out=116;              //668288-668319
                32'b0000000000001010001100101010xxxx: _out=116;              //668320-668335
                32'b00000000000010100011001010110xxx: _out=116;              //668336-668343
                
                32'b00000000000010100011001010111xxx: _out=117;              //668344-668351
                32'b00000000000010100011001011xxxxxx: _out=117;              //668352-668415
                32'b000000000000101000110011xxxxxxxx: _out=117;              //668416-668671
                32'b0000000000001010001101xxxxxxxxxx: _out=117;              //668672-669695
                32'b000000000000101000111xxxxxxxxxxx: _out=117;              //669696-671743
                32'b000000000000101001xxxxxxxxxxxxxx: _out=117;              //671744-688127
                32'b00000000000010101xxxxxxxxxxxxxxx: _out=117;              //688128-720895
                32'b000000000000101100xxxxxxxxxxxxxx: _out=117;              //720896-737279
                32'b0000000000001011010xxxxxxxxxxxxx: _out=117;              //737280-745471
                32'b00000000000010110110xxxxxxxxxxxx: _out=117;              //745472-749567
                32'b000000000000101101110000xxxxxxxx: _out=117;              //749568-749823
                32'b00000000000010110111000100xxxxxx: _out=117;              //749824-749887
                32'b000000000000101101110001010000xx: _out=117;              //749888-749891
                32'b0000000000001011011100010100010x: _out=117;              //749892-749893
                32'b00000000000010110111000101000110: _out=117;              //749894
                
                32'b00000000000010110111000101000111: _out=118;              //749895
                32'b00000000000010110111000101001xxx: _out=118;              //749896-749903
                32'b0000000000001011011100010101xxxx: _out=118;              //749904-749919
                32'b000000000000101101110001011xxxxx: _out=118;              //749920-749951
                32'b0000000000001011011100011xxxxxxx: _out=118;              //749952-750079
                32'b00000000000010110111001xxxxxxxxx: _out=118;              //750080-750591
                32'b0000000000001011011101xxxxxxxxxx: _out=118;              //750592-751615
                32'b000000000000101101111xxxxxxxxxxx: _out=118;              //751616-753663
                32'b00000000000010111xxxxxxxxxxxxxxx: _out=118;              //753664-786431
                32'b00000000000011000xxxxxxxxxxxxxxx: _out=118;              //786432-819199
                32'b000000000000110010xxxxxxxxxxxxxx: _out=118;              //819200-835583
                32'b00000000000011001100xxxxxxxxxxxx: _out=118;              //835584-839679
                32'b0000000000001100110100xxxxxxxxxx: _out=118;              //839680-840703
                32'b00000000000011001101010xxxxxxxxx: _out=118;              //840704-841215
                32'b0000000000001100110101100xxxxxxx: _out=118;              //841216-841343
                32'b000000000000110011010110100xxxxx: _out=118;              //841344-841375
                32'b0000000000001100110101101010xxxx: _out=118;              //841376-841391
                32'b000000000000110011010110101100xx: _out=118;              //841392-841395
                
                32'b000000000000110011010110101101xx: _out=119;              //841396-841399
                32'b00000000000011001101011010111xxx: _out=119;              //841400-841407
                32'b00000000000011001101011011xxxxxx: _out=119;              //841408-841471
                32'b000000000000110011010111xxxxxxxx: _out=119;              //841472-841727
                32'b000000000000110011011xxxxxxxxxxx: _out=119;              //841728-843775
                32'b0000000000001100111xxxxxxxxxxxxx: _out=119;              //843776-851967
                32'b0000000000001101xxxxxxxxxxxxxxxx: _out=119;              //851968-917503
                32'b000000000000111000xxxxxxxxxxxxxx: _out=119;              //917504-933887
                32'b0000000000001110010xxxxxxxxxxxxx: _out=119;              //933888-942079
                32'b0000000000001110011000xxxxxxxxxx: _out=119;              //942080-943103
                32'b00000000000011100110010xxxxxxxxx: _out=119;              //943104-943615
                32'b000000000000111001100110xxxxxxxx: _out=119;              //943616-943871
                32'b0000000000001110011001110xxxxxxx: _out=119;              //943872-943999
                32'b000000000000111001100111100xxxxx: _out=119;              //944000-944031
                32'b0000000000001110011001111010xxxx: _out=119;              //944032-944047
                32'b00000000000011100110011110110xxx: _out=119;              //944048-944055
                32'b000000000000111001100111101110xx: _out=119;              //944056-944059
                32'b00000000000011100110011110111100: _out=119;              //944060
                
                32'b00000000000011100110011110111101: _out=120;              //944061
                32'b0000000000001110011001111011111x: _out=120;              //944062-944063
                32'b00000000000011100110011111xxxxxx: _out=120;              //944064-944127
                32'b000000000000111001101xxxxxxxxxxx: _out=120;              //944128-946175
                32'b00000000000011100111xxxxxxxxxxxx: _out=120;              //946176-950271
                32'b00000000000011101xxxxxxxxxxxxxxx: _out=120;              //950272-983039
                32'b0000000000001111xxxxxxxxxxxxxxxx: _out=120;              //983040-1048575
                32'b0000000000010000000xxxxxxxxxxxxx: _out=120;              //1048576-1056767
                32'b000000000001000000100xxxxxxxxxxx: _out=120;              //1056768-1058815
                32'b000000000001000000101000xxxxxxxx: _out=120;              //1058816-1059071
                32'b0000000000010000001010010xxxxxxx: _out=120;              //1059072-1059199
                32'b000000000001000000101001100xxxxx: _out=120;              //1059200-1059231
                32'b0000000000010000001010011010xxxx: _out=120;              //1059232-1059247
                32'b000000000001000000101001101100xx: _out=120;              //1059248-1059251
                32'b0000000000010000001010011011010x: _out=120;              //1059252-1059253
                
                32'b0000000000010000001010011011011x: _out=121;              //1059254-1059255
                32'b00000000000100000010100110111xxx: _out=121;              //1059256-1059263
                32'b00000000000100000010100111xxxxxx: _out=121;              //1059264-1059327
                32'b00000000000100000010101xxxxxxxxx: _out=121;              //1059328-1059839
                32'b0000000000010000001011xxxxxxxxxx: _out=121;              //1059840-1060863
                32'b00000000000100000011xxxxxxxxxxxx: _out=121;              //1060864-1064959
                32'b000000000001000001xxxxxxxxxxxxxx: _out=121;              //1064960-1081343
                32'b00000000000100001xxxxxxxxxxxxxxx: _out=121;              //1081344-1114111
                32'b0000000000010001xxxxxxxxxxxxxxxx: _out=121;              //1114112-1179647
                32'b0000000000010010000xxxxxxxxxxxxx: _out=121;              //1179648-1187839
                32'b00000000000100100010000xxxxxxxxx: _out=121;              //1187840-1188351
                32'b0000000000010010001000100xxxxxxx: _out=121;              //1188352-1188479
                32'b0000000000010010001000101000xxxx: _out=121;              //1188480-1188495
                32'b000000000001001000100010100100xx: _out=121;              //1188496-1188499
                32'b0000000000010010001000101001010x: _out=121;              //1188500-1188501
                32'b00000000000100100010001010010110: _out=121;              //1188502
                
                32'b00000000000100100010001010010111: _out=122;              //1188503
                32'b00000000000100100010001010011xxx: _out=122;              //1188504-1188511
                32'b000000000001001000100010101xxxxx: _out=122;              //1188512-1188543
                32'b00000000000100100010001011xxxxxx: _out=122;              //1188544-1188607
                32'b000000000001001000100011xxxxxxxx: _out=122;              //1188608-1188863
                32'b0000000000010010001001xxxxxxxxxx: _out=122;              //1188864-1189887
                32'b000000000001001000101xxxxxxxxxxx: _out=122;              //1189888-1191935
                32'b00000000000100100011xxxxxxxxxxxx: _out=122;              //1191936-1196031
                32'b000000000001001001xxxxxxxxxxxxxx: _out=122;              //1196032-1212415
                32'b00000000000100101xxxxxxxxxxxxxxx: _out=122;              //1212416-1245183
                32'b0000000000010011xxxxxxxxxxxxxxxx: _out=122;              //1245184-1310719
                32'b000000000001010000xxxxxxxxxxxxxx: _out=122;              //1310720-1327103
                32'b00000000000101000100xxxxxxxxxxxx: _out=122;              //1327104-1331199
                32'b000000000001010001010xxxxxxxxxxx: _out=122;              //1331200-1333247
                32'b000000000001010001011000xxxxxxxx: _out=122;              //1333248-1333503
                32'b0000000000010100010110010000xxxx: _out=122;              //1333504-1333519
                32'b0000000000010100010110010001000x: _out=122;              //1333520-1333521
                
                32'b0000000000010100010110010001001x: _out=123;              //1333522-1333523
                32'b000000000001010001011001000101xx: _out=123;              //1333524-1333527
                32'b00000000000101000101100100011xxx: _out=123;              //1333528-1333535
                32'b000000000001010001011001001xxxxx: _out=123;              //1333536-1333567
                32'b00000000000101000101100101xxxxxx: _out=123;              //1333568-1333631
                32'b0000000000010100010110011xxxxxxx: _out=123;              //1333632-1333759
                32'b00000000000101000101101xxxxxxxxx: _out=123;              //1333760-1334271
                32'b0000000000010100010111xxxxxxxxxx: _out=123;              //1334272-1335295
                32'b0000000000010100011xxxxxxxxxxxxx: _out=123;              //1335296-1343487
                32'b00000000000101001xxxxxxxxxxxxxxx: _out=123;              //1343488-1376255
                32'b0000000000010101xxxxxxxxxxxxxxxx: _out=123;              //1376256-1441791
                32'b00000000000101100xxxxxxxxxxxxxxx: _out=123;              //1441792-1474559
                32'b000000000001011010xxxxxxxxxxxxxx: _out=123;              //1474560-1490943
                32'b00000000000101101100xxxxxxxxxxxx: _out=123;              //1490944-1495039
                32'b0000000000010110110100xxxxxxxxxx: _out=123;              //1495040-1496063
                32'b0000000000010110110101000xxxxxxx: _out=123;              //1496064-1496191
                32'b000000000001011011010100100xxxxx: _out=123;              //1496192-1496223
                32'b00000000000101101101010010100xxx: _out=123;              //1496224-1496231
                32'b000000000001011011010100101010xx: _out=123;              //1496232-1496235
                
                32'b000000000001011011010100101011xx: _out=124;              //1496236-1496239
                32'b0000000000010110110101001011xxxx: _out=124;              //1496240-1496255
                32'b00000000000101101101010011xxxxxx: _out=124;              //1496256-1496319
                32'b000000000001011011010101xxxxxxxx: _out=124;              //1496320-1496575
                32'b00000000000101101101011xxxxxxxxx: _out=124;              //1496576-1497087
                32'b000000000001011011011xxxxxxxxxxx: _out=124;              //1497088-1499135
                32'b0000000000010110111xxxxxxxxxxxxx: _out=124;              //1499136-1507327
                32'b0000000000010111xxxxxxxxxxxxxxxx: _out=124;              //1507328-1572863
                32'b0000000000011000xxxxxxxxxxxxxxxx: _out=124;              //1572864-1638399
                32'b00000000000110010xxxxxxxxxxxxxxx: _out=124;              //1638400-1671167
                32'b00000000000110011000xxxxxxxxxxxx: _out=124;              //1671168-1675263
                32'b000000000001100110010xxxxxxxxxxx: _out=124;              //1675264-1677311
                32'b0000000000011001100110xxxxxxxxxx: _out=124;              //1677312-1678335
                32'b000000000001100110011100xxxxxxxx: _out=124;              //1678336-1678591
                32'b0000000000011001100111010xxxxxxx: _out=124;              //1678592-1678719
                32'b00000000000110011001110110xxxxxx: _out=124;              //1678720-1678783
                32'b1100110011100000000000011100xxxx: _out=124;              //1678784-1678799
                32'b000000000001100110011101110100xx: _out=124;              //1678800-1678803
                32'b00000000000110011001110111010100: _out=124;              //1678804
                
                32'b00000000000110011001110111010101: _out=125;              //1678805
                32'b0000000000011001100111011101011x: _out=125;              //1678806-1678807
                32'b00000000000110011001110111011xxx: _out=125;              //1678808-1678815
                32'b000000000001100110011101111xxxxx: _out=125;              //1678816-1678847
                32'b00000000000110011001111xxxxxxxxx: _out=125;              //1678848-1679359
                32'b0000000000011001101xxxxxxxxxxxxx: _out=125;              //1679360-1687551
                32'b000000000001100111xxxxxxxxxxxxxx: _out=125;              //1687552-1703935
                32'b000000000001101xxxxxxxxxxxxxxxxx: _out=125;              //1703936-1835007
                32'b00000000000111000xxxxxxxxxxxxxxx: _out=125;              //1835008-1867775
                32'b0000000000011100100xxxxxxxxxxxxx: _out=125;              //1867776-1875967
                32'b00000000000111001010xxxxxxxxxxxx: _out=125;              //1875968-1880063
                32'b000000000001110010110xxxxxxxxxxx: _out=125;              //1880064-1882111
                32'b0000000000011100101110xxxxxxxxxx: _out=125;              //1882112-1883135
                32'b00000000000111001011110xxxxxxxxx: _out=125;              //1883136-1883647
                32'b0000000000011100101111100000000x: _out=125;              //1883648-1883649
                
                32'b0000000000011100101111100000001x: _out=126;              //1883650-1883651
                32'b000000000001110010111110000001xx: _out=126;              //1883652-1883655
                32'b00000000000111001011111000001xxx: _out=126;              //1883656-1883663
                32'b0000000000011100101111100001xxxx: _out=126;              //1883664-1883679
                32'b000000000001110010111110001xxxxx: _out=126;              //1883680-1883711
                32'b00000000000111001011111001xxxxxx: _out=126;              //1883712-1883775
                32'b0000000000011100101111101xxxxxxx: _out=126;              //1883776-1883903
                32'b000000000001110010111111xxxxxxxx: _out=126;              //1883904-1884159
                32'b000000000001110011xxxxxxxxxxxxxx: _out=126;              //1884160-1900543
                32'b0000000000011101xxxxxxxxxxxxxxxx: _out=126;              //1900544-1966079
                32'b000000000001111xxxxxxxxxxxxxxxxx: _out=126;              //1966080-2097151
                32'b0000000000100000000xxxxxxxxxxxxx: _out=126;              //2097152-2105343
                32'b00000000001000000010xxxxxxxxxxxx: _out=126;              //2105344-2109439
                32'b000000000010000000110xxxxxxxxxxx: _out=126;              //2109440-2111487
                32'b0000000000100000001110xxxxxxxxxx: _out=126;              //2111488-2112511
                32'b00000000001000000011110xxxxxxxxx: _out=126;              //2112512-2113023
                32'b000000000010000000111110xxxxxxxx: _out=126;              //2113024-2113279
                32'b0000000000100000001111110xxxxxxx: _out=126;              //2113280-2113407
                32'b00000000001000000011111110xxxxxx: _out=126;              //2113408-2113471
                32'b0000000000100000001111111100xxxx: _out=126;              //2113472-2113487
                32'b0000000000100000001111111101000x: _out=126;              //2113488-2113489
                
                32'b0000000000100000001111111101001x: _out=127;              //2113490-2113491
                32'b000000000010000000111111110101xx: _out=127;              //2113492-2113495
                32'b00000000001000000011111111011xxx: _out=127;              //2113496-2113503
                32'b000000000010000000111111111xxxxx: _out=127;              //2113504-2113535
                32'b000000000010000001xxxxxxxxxxxxxx: _out=127;              //2113536-2129919
                32'b00000000001000001xxxxxxxxxxxxxxx: _out=127;              //2129920-2162687
                32'b0000000000100001xxxxxxxxxxxxxxxx: _out=127;              //2162688-2228223
                32'b000000000010001xxxxxxxxxxxxxxxxx: _out=127;              //2228224-2359295
                32'b0000000000100100000xxxxxxxxxxxxx: _out=127;              //2359296-2367487
                32'b000000000010010000100xxxxxxxxxxx: _out=127;              //2367488-2369535
                32'b0000000000100100001010xxxxxxxxxx: _out=127;              //2369536-2370559
                32'b00000000001001000010110xxxxxxxxx: _out=127;              //2370560-2371071
                32'b000000000010010000101110xxxxxxxx: _out=127;              //2371072-2371327
                32'b000000000010010000101111000xxxxx: _out=127;              //2371328-2371359
                32'b00000000001001000010111100100xxx: _out=127;              //2371360-2371367
                32'b000000000010010000101111001010xx: _out=127;              //2371368-2371371
                32'b0000000000100100001011110010110x: _out=127;              //2371372-2371373
                
                32'b0000000000100100001011110010111x: _out=128;              //2371374-2371375
                32'b0000000000100100001011110011xxxx: _out=128;              //2371376-2371391
                32'b00000000001001000010111101xxxxxx: _out=128;              //2371392-2371455
                32'b0000000000100100001011111xxxxxxx: _out=128;              //2371456-2371583
                32'b00000000001001000011xxxxxxxxxxxx: _out=128;              //2371584-2375679
                32'b000000000010010001xxxxxxxxxxxxxx: _out=128;              //2375680-2392063
                32'b00000000001001001xxxxxxxxxxxxxxx: _out=128;              //2392064-2424831
                32'b0000000000100101xxxxxxxxxxxxxxxx: _out=128;              //2424832-2490367
                32'b000000000010011xxxxxxxxxxxxxxxxx: _out=128;              //2490368-2621439
                32'b00000000001010000xxxxxxxxxxxxxxx: _out=128;              //2621440-2654207
                32'b00000000001010001000xxxxxxxxxxxx: _out=128;              //2654208-2658303
                32'b000000000010100010010xxxxxxxxxxx: _out=128;              //2658304-2660351
                32'b000000000010100010011000xxxxxxxx: _out=128;              //2660352-2660607
                32'b00000000001010001001100100xxxxxx: _out=128;              //2660608-2660671
                32'b000000000010100010011001010xxxxx: _out=128;              //2660672-2660703
                32'b0000000000101000100110010110xxxx: _out=128;              //2660704-2660719
                32'b000000000010100010011001011100xx: _out=128;              //2660720-2660723
                32'b0000000000101000100110010111010x: _out=128;              //2660724-2660725
                
                32'b0000000000101000100110010111011x: _out=129;              //2660726-2660727
                32'b00000000001010001001100101111xxx: _out=129;              //2660728-2660735
                32'b0000000000101000100110011xxxxxxx: _out=129;              //2660736-2660863
                32'b00000000001010001001101xxxxxxxxx: _out=129;              //2660864-2661375
                32'b0000000000101000100111xxxxxxxxxx: _out=129;              //2661376-2662399
                32'b0000000000101000101xxxxxxxxxxxxx: _out=129;              //2662400-2670591
                32'b000000000010100011xxxxxxxxxxxxxx: _out=129;              //2670592-2686975
                32'b0000000000101001xxxxxxxxxxxxxxxx: _out=129;              //2686976-2752511
                32'b000000000010101xxxxxxxxxxxxxxxxx: _out=129;              //2752512-2883583
                32'b0000000000101100xxxxxxxxxxxxxxxx: _out=129;              //2883584-2949119
                32'b00000000001011010xxxxxxxxxxxxxxx: _out=129;              //2949120-2981887
                32'b000000000010110110000xxxxxxxxxxx: _out=129;              //2981888-2983935
                32'b0000000000101101100010xxxxxxxxxx: _out=129;              //2983936-2984959
                32'b000000000010110110001100xxxxxxxx: _out=129;              //2984960-2985215
                32'b0000000000101101100011010xxxxxxx: _out=129;              //2985216-2985343
                32'b000000000010110110001101100xxxxx: _out=129;              //2985344-2985375
                32'b000000000010110110001101101000xx: _out=129;              //2985376-2985379
                32'b0000000000101101100011011010010x: _out=129;              //2985380-2985381
                32'b00000000001011011000110110100110: _out=129;              //2985382
                
                32'b00000000001011011000110110100111: _out=130;              //2985383
                32'b00000000001011011000110110101xxx: _out=130;              //2985384-2985391
                32'b0000000000101101100011011011xxxx: _out=130;              //2985392-2985407
                32'b00000000001011011000110111xxxxxx: _out=130;              //2985408-2985471
                32'b00000000001011011000111xxxxxxxxx: _out=130;              //2985472-2985983
                32'b00000000001011011001xxxxxxxxxxxx: _out=130;              //2985984-2990079
                32'b0000000000101101101xxxxxxxxxxxxx: _out=130;              //2990080-2998271
                32'b000000000010110111xxxxxxxxxxxxxx: _out=130;              //2998272-3014655
                32'b000000000010111xxxxxxxxxxxxxxxxx: _out=130;              //3014656-3145727
                32'b000000000011000xxxxxxxxxxxxxxxxx: _out=130;              //3145728-3276799
                32'b0000000000110010xxxxxxxxxxxxxxxx: _out=130;              //3276800-3342335
                32'b00000000001100110000xxxxxxxxxxxx: _out=130;              //3342336-3346431
                32'b000000000011001100010xxxxxxxxxxx: _out=130;              //3346432-3348479
                32'b0000000000110011000110xxxxxxxxxx: _out=130;              //3348480-3349503
                32'b0000000000110011000111000xxxxxxx: _out=130;              //3349504-3349631
                32'b0000000000110011000111001000xxxx: _out=130;              //3349632-3349647
                32'b000000000011001100011100100100xx: _out=130;              //3349648-3349651
                32'b0000000000110011000111001001010x: _out=130;              //3349652-3349653
                32'b00000000001100110001110010010110: _out=130;              //3349654
                
                32'b00000000001100110001110010010111: _out=131;              //3349655
                32'b00000000001100110001110010011xxx: _out=131;              //3349656-3349663
                32'b000000000011001100011100101xxxxx: _out=131;              //3349664-3349695
                32'b00000000001100110001110011xxxxxx: _out=131;              //3349696-3349759
                32'b000000000011001100011101xxxxxxxx: _out=131;              //3349760-3350015
                32'b00000000001100110001111xxxxxxxxx: _out=131;              //3350016-3350527
                32'b0000000000110011001xxxxxxxxxxxxx: _out=131;              //3350528-3358719
                32'b000000000011001101xxxxxxxxxxxxxx: _out=131;              //3358720-3375103
                32'b00000000001100111xxxxxxxxxxxxxxx: _out=131;              //3375104-3407871
                32'b00000000001101xxxxxxxxxxxxxxxxxx: _out=131;              //3407872-3670015
                32'b0000000000111000xxxxxxxxxxxxxxxx: _out=131;              //3670016-3735551
                32'b000000000011100100xxxxxxxxxxxxxx: _out=131;              //3735552-3751935
                32'b00000000001110010100xxxxxxxxxxxx: _out=131;              //3751936-3756031
                32'b000000000011100101010xxxxxxxxxxx: _out=131;              //3756032-3758079
                32'b000000000011100101011000xxxxxxxx: _out=131;              //3758080-3758335
                32'b000000000011100101011001000xxxxx: _out=131;              //3758336-3758367
                32'b000000000011100101011001001000xx: _out=131;              //3758368-3758371
                32'b0000000000111001010110010010010x: _out=131;              //3758372-3758373
                32'b00000000001110010101100100100110: _out=131;              //3758374
                
                32'b00000000001110010101100100100111: _out=132;              //3758375
                32'b00000000001110010101100100101xxx: _out=132;              //3758376-3758383
                32'b0000000000111001010110010011xxxx: _out=132;              //3758384-3758399
                32'b00000000001110010101100101xxxxxx: _out=132;              //3758400-3758463
                32'b0000000000111001010110011xxxxxxx: _out=132;              //3758464-3758591
                32'b00000000001110010101101xxxxxxxxx: _out=132;              //3758592-3759103
                32'b0000000000111001010111xxxxxxxxxx: _out=132;              //3759104-3760127
                32'b0000000000111001011xxxxxxxxxxxxx: _out=132;              //3760128-3768319
                32'b00000000001110011xxxxxxxxxxxxxxx: _out=132;              //3768320-3801087
                32'b000000000011101xxxxxxxxxxxxxxxxx: _out=132;              //3801088-3932159
                32'b00000000001111xxxxxxxxxxxxxxxxxx: _out=132;              //3932160-4194303
                32'b000000000100000000xxxxxxxxxxxxxx: _out=132;              //4194304-4210687
                32'b00000000010000000100xxxxxxxxxxxx: _out=132;              //4210688-4214783
                32'b000000000100000001010xxxxxxxxxxx: _out=132;              //4214784-4216831
                32'b0000000001000000010110000xxxxxxx: _out=132;              //4216832-4216959
                32'b000000000100000001011000100000xx: _out=132;              //4216960-4216963
                32'b0000000001000000010110001000010x: _out=132;              //4216964-4216965
                
                32'b0000000001000000010110001000011x: _out=133;              //4216966-4216967
                32'b00000000010000000101100010001xxx: _out=133;              //4216968-4216975
                32'b0000000001000000010110001001xxxx: _out=133;              //4216976-4216991
                32'b000000000100000001011000101xxxxx: _out=133;              //4216992-4217023
                32'b00000000010000000101100011xxxxxx: _out=133;              //4217024-4217087
                32'b000000000100000001011001xxxxxxxx: _out=133;              //4217088-4217343
                32'b00000000010000000101101xxxxxxxxx: _out=133;              //4217344-4217855
                32'b0000000001000000010111xxxxxxxxxx: _out=133;              //4217856-4218879
                32'b0000000001000000011xxxxxxxxxxxxx: _out=133;              //4218880-4227071
                32'b00000000010000001xxxxxxxxxxxxxxx: _out=133;              //4227072-4259839
                32'b0000000001000001xxxxxxxxxxxxxxxx: _out=133;              //4259840-4325375
                32'b000000000100001xxxxxxxxxxxxxxxxx: _out=133;              //4325376-4456447
                32'b00000000010001xxxxxxxxxxxxxxxxxx: _out=133;              //4456448-4718591
                32'b0000000001001000000xxxxxxxxxxxxx: _out=133;              //4718592-4726783
                32'b00000000010010000010xxxxxxxxxxxx: _out=133;              //4726784-4730879
                32'b00000000010010000011000xxxxxxxxx: _out=133;              //4730880-4731391
                32'b00000000010010000011001000xxxxxx: _out=133;              //4731392-4731455
                32'b000000000100100000110010010xxxxx: _out=133;              //4731456-4731487
                32'b0000000001001000001100100110xxxx: _out=133;              //4731488-4731503
                32'b00000000010010000011001001110xxx: _out=133;              //4731504-4731511
                32'b00000000010010000011001001111000: _out=133;              //4731512
                
                32'b00000000010010000011001001111001: _out=134;              //4731513
                32'b0000000001001000001100100111101x: _out=134;              //4731514-4731515
                32'b000000000100100000110010011111xx: _out=134;              //4731516-4731519
                32'b0000000001001000001100101xxxxxxx: _out=134;              //4731520-4731647
                32'b000000000100100000110011xxxxxxxx: _out=134;              //4731648-4731903
                32'b0000000001001000001101xxxxxxxxxx: _out=134;              //4731904-4732927
                32'b000000000100100000111xxxxxxxxxxx: _out=134;              //4732928-4734975
                32'b000000000100100001xxxxxxxxxxxxxx: _out=134;              //4734976-4751359
                32'b00000000010010001xxxxxxxxxxxxxxx: _out=134;              //4751360-4784127
                32'b0000000001001001xxxxxxxxxxxxxxxx: _out=134;              //4784128-4849663
                32'b000000000100101xxxxxxxxxxxxxxxxx: _out=134;              //4849664-4980735
                32'b00000000010011xxxxxxxxxxxxxxxxxx: _out=134;              //4980736-5242879
                32'b0000000001010000xxxxxxxxxxxxxxxx: _out=134;              //5242880-5308415
                32'b000000000101000100000000xxxxxxxx: _out=134;              //5308416-5308671
                32'b0000000001010001000000010xxxxxxx: _out=134;              //5308672-5308799
                32'b000000000101000100000001100xxxxx: _out=134;              //5308800-5308831
                32'b00000000010100010000000110100xxx: _out=134;              //5308832-5308839
                32'b000000000101000100000001101010xx: _out=134;              //5308840-5308843
                32'b00000000010100010000000110101100: _out=134;              //5308844
                
                32'b00000000010100010000000110101101: _out=135;              //5308845
                32'b0000000001010001000000011010111x: _out=135;              //5308846-5308847
                32'b0000000001010001000000011011xxxx: _out=135;              //5308848-5308863
                32'b00000000010100010000000111xxxxxx: _out=135;              //5308864-5308927
                32'b00000000010100010000001xxxxxxxxx: _out=135;              //5308928-5309439
                32'b0000000001010001000001xxxxxxxxxx: _out=135;              //5309440-5310463
                32'b000000000101000100001xxxxxxxxxxx: _out=135;              //5310464-5312511
                32'b00000000010100010001xxxxxxxxxxxx: _out=135;              //5312512-5316607
                32'b0000000001010001001xxxxxxxxxxxxx: _out=135;              //5316608-5324799
                32'b000000000101000101xxxxxxxxxxxxxx: _out=135;              //5324800-5341183
                32'b00000000010100011xxxxxxxxxxxxxxx: _out=135;              //5341184-5373951
                32'b000000000101001xxxxxxxxxxxxxxxxx: _out=135;              //5373952-5505023
                32'b00000000010101xxxxxxxxxxxxxxxxxx: _out=135;              //5505024-5767167
                32'b000000000101100xxxxxxxxxxxxxxxxx: _out=135;              //5767168-5898239
                32'b00000000010110100xxxxxxxxxxxxxxx: _out=135;              //5898240-5931007
                32'b000000000101101010xxxxxxxxxxxxxx: _out=135;              //5931008-5947391
                32'b0000000001011010110xxxxxxxxxxxxx: _out=135;              //5947392-5955583
                32'b0000000001011010111000xxxxxxxxxx: _out=135;              //5955584-5956607
                32'b00000000010110101110010000000xxx: _out=135;              //5956608-5956615
                32'b000000000101101011100100000010xx: _out=135;              //5956616-5956619
                32'b0000000001011010111001000000110x: _out=135;              //5956620-5956621
                
                32'b0000000001011010111001000000111x: _out=136;              //5956622-5956623
                32'b0000000001011010111001000001xxxx: _out=136;              //5956624-5956639
                32'b000000000101101011100100001xxxxx: _out=136;              //5956640-5956671
                32'b00000000010110101110010001xxxxxx: _out=136;              //5956672-5956735
                32'b0000000001011010111001001xxxxxxx: _out=136;              //5956736-5956863
                32'b000000000101101011100101xxxxxxxx: _out=136;              //5956864-5957119
                32'b00000000010110101110011xxxxxxxxx: _out=136;              //5957120-5957631
                32'b000000000101101011101xxxxxxxxxxx: _out=136;              //5957632-5959679
                32'b00000000010110101111xxxxxxxxxxxx: _out=136;              //5959680-5963775
                32'b0000000001011011xxxxxxxxxxxxxxxx: _out=136;              //5963776-6029311
                32'b00000000010111xxxxxxxxxxxxxxxxxx: _out=136;              //6029312-6291455
                32'b00000000011000xxxxxxxxxxxxxxxxxx: _out=136;              //6291456-6553599
                32'b0000000001100100xxxxxxxxxxxxxxxx: _out=136;              //6553600-6619135
                32'b00000000011001010xxxxxxxxxxxxxxx: _out=136;              //6619136-6651903
                32'b000000000110010110xxxxxxxxxxxxxx: _out=136;              //6651904-6668287
                32'b0000000001100101110xxxxxxxxxxxxx: _out=136;              //6668288-6676479
                32'b00000000011001011110xxxxxxxxxxxx: _out=136;              //6676480-6680575
                32'b000000000110010111110xxxxxxxxxxx: _out=136;              //6680576-6682623
                32'b00000000011001011111100xxxxxxxxx: _out=136;              //6682624-6683135
                32'b000000000110010111111010xxxxxxxx: _out=136;              //6683136-6683391
                32'b000000000110010111111011000xxxxx: _out=136;              //6683392-6683423
                32'b0000000001100101111110110010xxxx: _out=136;              //6683424-6683439
                
                32'b0000000001100101111110110011xxxx: _out=137;              //6683440-6683455
                32'b00000000011001011111101101xxxxxx: _out=137;              //6683456-6683519
                32'b0000000001100101111110111xxxxxxx: _out=137;              //6683520-6683647
                32'b0000000001100101111111xxxxxxxxxx: _out=137;              //6683648-6684671
                32'b000000000110011xxxxxxxxxxxxxxxxx: _out=137;              //6684672-6815743
                32'b0000000001101xxxxxxxxxxxxxxxxxxx: _out=137;              //6815744-7340031
                32'b000000000111000xxxxxxxxxxxxxxxxx: _out=137;              //7340032-7471103
                32'b000000000111001000xxxxxxxxxxxxxx: _out=137;              //7471104-7487487
                32'b0000000001110010010xxxxxxxxxxxxx: _out=137;              //7487488-7495679
                32'b000000000111001001100xxxxxxxxxxx: _out=137;              //7495680-7497727
                32'b0000000001110010011010xxxxxxxxxx: _out=137;              //7497728-7498751
                32'b0000000001110010011011000xxxxxxx: _out=137;              //7498752-7498879
                32'b000000000111001001101100100xxxxx: _out=137;              //7498880-7498911
                32'b0000000001110010011011001010xxxx: _out=137;              //7498912-7498927
                32'b00000000011100100110110010110xxx: _out=137;              //7498928-7498935
                32'b000000000111001001101100101110xx: _out=137;              //7498936-7498939
                32'b0000000001110010011011001011110x: _out=137;              //7498940-7498941
                32'b00000000011100100110110010111110: _out=137;              //7498942
                
                32'b00000000011100100110110010111111: _out=138;              //7498943
                32'b00000000011100100110110011xxxxxx: _out=138;              //7498944-7499007
                32'b000000000111001001101101xxxxxxxx: _out=138;              //7499008-7499263
                32'b00000000011100100110111xxxxxxxxx: _out=138;              //7499264-7499775
                32'b00000000011100100111xxxxxxxxxxxx: _out=138;              //7499776-7503871
                32'b00000000011100101xxxxxxxxxxxxxxx: _out=138;              //7503872-7536639
                32'b0000000001110011xxxxxxxxxxxxxxxx: _out=138;              //7536640-7602175
                32'b00000000011101xxxxxxxxxxxxxxxxxx: _out=138;              //7602176-7864319
                32'b0000000001111xxxxxxxxxxxxxxxxxxx: _out=138;              //7864320-8388607
                32'b000000001000000000xxxxxxxxxxxxxx: _out=138;              //8388608-8404991
                32'b0000000010000000010xxxxxxxxxxxxx: _out=138;              //8404992-8413183
                32'b00000000100000000110000xxxxxxxxx: _out=138;              //8413184-8413695
                32'b000000001000000001100010xxxxxxxx: _out=138;              //8413696-8413951
                
                32'b000000001000000001100011xxxxxxxx: _out=139;              //8413952-8414207
                32'b0000000010000000011001xxxxxxxxxx: _out=139;              //8414208-8415231
                32'b000000001000000001101xxxxxxxxxxx: _out=139;              //8415232-8417279
                32'b00000000100000000111xxxxxxxxxxxx: _out=139;              //8417280-8421375
                32'b00000000100000001xxxxxxxxxxxxxxx: _out=139;              //8421376-8454143
                32'b0000000010000001xxxxxxxxxxxxxxxx: _out=139;              //8454144-8519679
                32'b000000001000001xxxxxxxxxxxxxxxxx: _out=139;              //8519680-8650751
                32'b00000000100001xxxxxxxxxxxxxxxxxx: _out=139;              //8650752-8912895
                32'b0000000010001xxxxxxxxxxxxxxxxxxx: _out=139;              //8912896-9437183
                32'b000000001001000000000xxxxxxxxxxx: _out=139;              //9437184-9439231
                32'b0000000010010000000010xxxxxxxxxx: _out=139;              //9439232-9440255
                32'b000000001001000000001100xxxxxxxx: _out=139;              //9440256-9440511
                32'b00000000100100000000110100xxxxxx: _out=139;              //9440512-9440575
                32'b000000001001000000001101010xxxxx: _out=139;              //9440576-9440607
                32'b00000000100100000000110101100000: _out=139;              //9440608
                
                32'b00000000100100000000110101100001: _out=140;              //9440609
                32'b0000000010010000000011010110001x: _out=140;              //9440610-9440611
                32'b000000001001000000001101011001xx: _out=140;              //9440612-9440615
                32'b00000000100100000000110101101xxx: _out=140;              //9440616-9440623
                32'b0000000010010000000011010111xxxx: _out=140;              //9440624-9440639
                32'b0000000010010000000011011xxxxxxx: _out=140;              //9440640-9440767
                32'b00000000100100000000111xxxxxxxxx: _out=140;              //9440768-9441279
                32'b00000000100100000001xxxxxxxxxxxx: _out=140;              //9441280-9445375
                32'b0000000010010000001xxxxxxxxxxxxx: _out=140;              //9445376-9453567
                32'b000000001001000001xxxxxxxxxxxxxx: _out=140;              //9453568-9469951
                32'b00000000100100001xxxxxxxxxxxxxxx: _out=140;              //9469952-9502719
                32'b0000000010010001xxxxxxxxxxxxxxxx: _out=140;              //9502720-9568255
                32'b000000001001001xxxxxxxxxxxxxxxxx: _out=140;              //9568256-9699327
                32'b00000000100101xxxxxxxxxxxxxxxxxx: _out=140;              //9699328-9961471
                32'b0000000010011xxxxxxxxxxxxxxxxxxx: _out=140;              //9961472-10485759
                32'b0000000010100000xxxxxxxxxxxxxxxx: _out=140;              //10485760-10551295
                32'b00000000101000010xxxxxxxxxxxxxxx: _out=140;              //10551296-10584063
                32'b0000000010100001100xxxxxxxxxxxxx: _out=140;              //10584064-10592255
                32'b000000001010000110100000xxxxxxxx: _out=140;              //10592256-10592511
                32'b0000000010100001101000010000xxxx: _out=140;              //10592512-10592527
                32'b00000000101000011010000100010xxx: _out=140;              //10592528-10592535
                32'b0000000010100001101000010001100x: _out=140;              //10592536-10592537

                32'b0000000010100001101000010001101x: _out=141;              //10592538-10592539
                32'b000000001010000110100001000111xx: _out=141;              //10592540-10592543
                32'b000000001010000110100001001xxxxx: _out=141;              //10592544-10592575
                32'b00000000101000011010000101xxxxxx: _out=141;              //10592576-10592639
                32'b0000000010100001101000011xxxxxxx: _out=141;              //10592640-10592767
                32'b00000000101000011010001xxxxxxxxx: _out=141;              //10592768-10593279
                32'b0000000010100001101001xxxxxxxxxx: _out=141;              //10593280-10594303
                32'b000000001010000110101xxxxxxxxxxx: _out=141;              //10594304-10596351
                32'b00000000101000011011xxxxxxxxxxxx: _out=141;              //10596352-10600447
                32'b000000001010000111xxxxxxxxxxxxxx: _out=141;              //10600448-10616831
                32'b000000001010001xxxxxxxxxxxxxxxxx: _out=141;              //10616832-10747903
                32'b00000000101001xxxxxxxxxxxxxxxxxx: _out=141;              //10747904-11010047
                32'b0000000010101xxxxxxxxxxxxxxxxxxx: _out=141;              //11010048-11534335
                32'b00000000101100xxxxxxxxxxxxxxxxxx: _out=141;              //11534336-11796479
                32'b0000000010110100xxxxxxxxxxxxxxxx: _out=141;              //11796480-11862015
                32'b000000001011010100xxxxxxxxxxxxxx: _out=141;              //11862016-11878399
                32'b00000000101101010100xxxxxxxxxxxx: _out=141;              //11878400-11882495
                32'b000000001011010101010xxxxxxxxxxx: _out=141;              //11882496-11884543
                32'b000000001011010101011000xxxxxxxx: _out=141;              //11884544-11884799
                32'b0000000010110101010110010xxxxxxx: _out=141;              //11884800-11884927
                32'b00000000101101010101100110xxxxxx: _out=141;              //11884928-11884991
                32'b0000000010110101010110011100xxxx: _out=141;              //11884992-11885007
                32'b00000000101101010101100111010xxx: _out=141;              //11885008-11885015
                32'b000000001011010101011001110110xx: _out=141;              //11885016-11885019
                32'b0000000010110101010110011101110x: _out=141;              //11885020-11885021
                32'b00000000101101010101100111011110: _out=141;              //11885022

                32'b00000000101101010101100111011111: _out=142;              //11885023
                32'b000000001011010101011001111xxxxx: _out=142;              //11885024-11885055
                32'b00000000101101010101101xxxxxxxxx: _out=142;              //11885056-11885567
                32'b0000000010110101010111xxxxxxxxxx: _out=142;              //11885568-11886591
                32'b0000000010110101011xxxxxxxxxxxxx: _out=142;              //11886592-11894783
                32'b00000000101101011xxxxxxxxxxxxxxx: _out=142;              //11894784-11927551
                32'b000000001011011xxxxxxxxxxxxxxxxx: _out=142;              //11927552-12058623
                32'b0000000010111xxxxxxxxxxxxxxxxxxx: _out=142;              //12058624-12582911
                32'b0000000011000xxxxxxxxxxxxxxxxxxx: _out=142;              //12582912-13107199
                32'b000000001100100xxxxxxxxxxxxxxxxx: _out=142;              //13107200-13238271
                32'b0000000011001010xxxxxxxxxxxxxxxx: _out=142;              //13238272-13303807
                32'b000000001100101100xxxxxxxxxxxxxx: _out=142;              //13303808-13320191
                32'b0000000011001011010xxxxxxxxxxxxx: _out=142;              //13320192-13328383
                32'b00000000110010110110xxxxxxxxxxxx: _out=142;              //13328384-13332479
                32'b000000001100101101110xxxxxxxxxxx: _out=142;              //13332480-13334527
                32'b00000000110010110111100xxxxxxxxx: _out=142;              //13334528-13335039
                32'b0000000011001011011110100xxxxxxx: _out=142;              //13335040-13335167
                32'b000000001100101101111010100xxxxx: _out=142;              //13335168-13335199
                32'b00000000110010110111101010100xxx: _out=142;              //13335200-13335207
                32'b000000001100101101111010101010xx: _out=142;              //13335208-13335211
                32'b0000000011001011011110101010110x: _out=142;              //13335212-13335213
                32'b00000000110010110111101010101110: _out=142;              //13335214
                
                32'b00000000110010110111101010101111: _out=143;              //13335215
                32'b0000000011001011011110101011xxxx: _out=143;              //13335216-13335231
                32'b00000000110010110111101011xxxxxx: _out=143;              //13335232-13335295
                32'b000000001100101101111011xxxxxxxx: _out=143;              //13335296-13335551
                32'b0000000011001011011111xxxxxxxxxx: _out=143;              //13335552-13336575
                32'b00000000110010111xxxxxxxxxxxxxxx: _out=143;              //13336576-13369343
                32'b00000000110011xxxxxxxxxxxxxxxxxx: _out=143;              //13369344-13631487
                32'b000000001101xxxxxxxxxxxxxxxxxxxx: _out=143;              //13631488-14680063
                32'b00000000111000xxxxxxxxxxxxxxxxxx: _out=143;              //14680064-14942207
                32'b000000001110010000xxxxxxxxxxxxxx: _out=143;              //14942208-14958591
                32'b000000001110010001000xxxxxxxxxxx: _out=143;              //14958592-14960639
                32'b0000000011100100010010xxxxxxxxxx: _out=143;              //14960640-14961663
                32'b00000000111001000100110xxxxxxxxx: _out=143;              //14961664-14962175
                32'b0000000011100100010011100xxxxxxx: _out=143;              //14962176-14962303
                32'b000000001110010001001110100xxxxx: _out=143;              //14962304-14962335
                32'b0000000011100100010011101010xxxx: _out=143;              //14962336-14962351
                32'b000000001110010001001110101100xx: _out=143;              //14962352-14962355
                32'b00000000111001000100111010110100: _out=143;              //14962356
                
                32'b00000000111001000100111010110101: _out=144;              //14962357
                32'b0000000011100100010011101011011x: _out=144;              //14962358-14962359
                32'b00000000111001000100111010111xxx: _out=144;              //14962360-14962367
                32'b00000000111001000100111011xxxxxx: _out=144;              //14962368-14962431
                32'b000000001110010001001111xxxxxxxx: _out=144;              //14962432-14962687
                32'b00000000111001000101xxxxxxxxxxxx: _out=144;              //14962688-14966783
                32'b0000000011100100011xxxxxxxxxxxxx: _out=144;              //14966784-14974975
                32'b00000000111001001xxxxxxxxxxxxxxx: _out=144;              //14974976-15007743
                32'b0000000011100101xxxxxxxxxxxxxxxx: _out=144;              //15007744-15073279
                32'b000000001110011xxxxxxxxxxxxxxxxx: _out=144;              //15073280-15204351
                32'b0000000011101xxxxxxxxxxxxxxxxxxx: _out=144;              //15204352-15728639
                32'b000000001111xxxxxxxxxxxxxxxxxxxx: _out=144;              //15728640-16777215
                32'b0000000100000000000xxxxxxxxxxxxx: _out=144;              //16777216-16785407
                32'b000000010000000000100xxxxxxxxxxx: _out=144;              //16785408-16787455
                32'b00000001000000000010100xxxxxxxxx: _out=144;              //16787456-16787967
                32'b00000001000000000010101000xxxxxx: _out=144;              //16787968-16788031
                32'b00000001000000000010101001000xxx: _out=144;              //16788032-16788039
                32'b00000001000000000010101001001000: _out=144;              //16788040
                
                32'b00000001000000000010101001001001: _out=145;              //16788041
                32'b0000000100000000001010100100101x: _out=145;              //16788042-16788043
                32'b000000010000000000101010010011xx: _out=145;              //16788044-16788047
                32'b0000000100000000001010100101xxxx: _out=145;              //16788048-16788063
                32'b000000010000000000101010011xxxxx: _out=145;              //16788064-16788095
                32'b0000000100000000001010101xxxxxxx: _out=145;              //16788096-16788223
                32'b000000010000000000101011xxxxxxxx: _out=145;              //16788224-16788479
                32'b0000000100000000001011xxxxxxxxxx: _out=145;              //16788480-16789503
                32'b00000001000000000011xxxxxxxxxxxx: _out=145;              //16789504-16793599
                32'b000000010000000001xxxxxxxxxxxxxx: _out=145;              //16793600-16809983
                32'b00000001000000001xxxxxxxxxxxxxxx: _out=145;              //16809984-16842751
                32'b0000000100000001xxxxxxxxxxxxxxxx: _out=145;              //16842752-16908287
                32'b000000010000001xxxxxxxxxxxxxxxxx: _out=145;              //16908288-17039359
                32'b00000001000001xxxxxxxxxxxxxxxxxx: _out=145;              //17039360-17301503
                32'b0000000100001xxxxxxxxxxxxxxxxxxx: _out=145;              //17301504-17825791
                32'b0000000100010xxxxxxxxxxxxxxxxxxx: _out=145;              //17825792-18350079
                32'b00000001000110xxxxxxxxxxxxxxxxxx: _out=145;              //18350080-18612223
                32'b000000010001110xxxxxxxxxxxxxxxxx: _out=145;              //18612224-18743295
                32'b0000000100011110xxxxxxxxxxxxxxxx: _out=145;              //18743296-18808831
                32'b000000010001111100xxxxxxxxxxxxxx: _out=145;              //18808832-18825215
                32'b0000000100011111010xxxxxxxxxxxxx: _out=145;              //18825216-18833407
                32'b000000010001111101100xxxxxxxxxxx: _out=145;              //18833408-18835455
                32'b0000000100011111011010xxxxxxxxxx: _out=145;              //18835456-18836479
                32'b00000001000111110110110000000xxx: _out=145;              //18836480-18836487
                32'b0000000100011111011011000000100x: _out=145;              //18836488-18836489
                32'b00000001000111110110110000001010: _out=145;              //18836490
                
                32'b00000001000111110110110000001011: _out=146;              //18836491
                32'b000000010001111101101100000011xx: _out=146;              //18836492-18836495
                32'b0000000100011111011011000001xxxx: _out=146;              //18836496-18836511
                32'b000000010001111101101100001xxxxx: _out=146;              //18836512-18836543
                32'b00000001000111110110110001xxxxxx: _out=146;              //18836544-18836607
                32'b0000000100011111011011001xxxxxxx: _out=146;              //18836608-18836735
                32'b000000010001111101101101xxxxxxxx: _out=146;              //18836736-18836991
                32'b00000001000111110110111xxxxxxxxx: _out=146;              //18836992-18837503
                32'b00000001000111110111xxxxxxxxxxxx: _out=146;              //18837504-18841599
                32'b00000001000111111xxxxxxxxxxxxxxx: _out=146;              //18841600-18874367
                32'b00000001001xxxxxxxxxxxxxxxxxxxxx: _out=146;              //18874368-20971519
                32'b000000010100000xxxxxxxxxxxxxxxxx: _out=146;              //20971520-21102591
                32'b000000010100001000xxxxxxxxxxxxxx: _out=146;              //21102592-21118975
                32'b0000000101000010010xxxxxxxxxxxxx: _out=146;              //21118976-21127167
                32'b00000001010000100110xxxxxxxxxxxx: _out=146;              //21127168-21131263
                32'b000000010100001001110xxxxxxxxxxx: _out=146;              //21131264-21133311
                32'b0000000101000010011110xxxxxxxxxx: _out=146;              //21133312-21134335
                32'b00000001010000100111110xxxxxxxxx: _out=146;              //21134336-21134847
                32'b000000010100001001111110000xxxxx: _out=146;              //21134848-21134879
                32'b00000001010000100111111000100xxx: _out=146;              //21134880-21134887
                32'b0000000101000010011111100010100x: _out=146;              //21134888-21134889
                32'b00000001010000100111111000101010: _out=146;              //21134890
                
                32'b00000001010000100111111000101011: _out=147;              //21134891
                32'b000000010100001001111110001011xx: _out=147;              //21134892-21134895
                32'b0000000101000010011111100011xxxx: _out=147;              //21134896-21134911
                32'b00000001010000100111111001xxxxxx: _out=147;              //21134912-21134975
                32'b0000000101000010011111101xxxxxxx: _out=147;              //21134976-21135103
                32'b000000010100001001111111xxxxxxxx: _out=147;              //21135104-21135359
                32'b00000001010000101xxxxxxxxxxxxxxx: _out=147;              //21135360-21168127
                32'b0000000101000011xxxxxxxxxxxxxxxx: _out=147;              //21168128-21233663
                32'b00000001010001xxxxxxxxxxxxxxxxxx: _out=147;              //21233664-21495807
                32'b0000000101001xxxxxxxxxxxxxxxxxxx: _out=147;              //21495808-22020095
                32'b000000010101xxxxxxxxxxxxxxxxxxxx: _out=147;              //22020096-23068671
                32'b0000000101100xxxxxxxxxxxxxxxxxxx: _out=147;              //23068672-23592959
                32'b0000000101101000xxxxxxxxxxxxxxxx: _out=147;              //23592960-23658495
                32'b00000001011010010xxxxxxxxxxxxxxx: _out=147;              //23658496-23691263
                32'b000000010110100110xxxxxxxxxxxxxx: _out=147;              //23691264-23707647
                32'b00000001011010011100xxxxxxxxxxxx: _out=147;              //23707648-23711743
                32'b0000000101101001110100xxxxxxxxxx: _out=147;              //23711744-23712767
                32'b00000001011010011101010xxxxxxxxx: _out=147;              //23712768-23713279
                32'b000000010110100111010110xxxxxxxx: _out=147;              //23713280-23713535
                32'b0000000101101001110101110xxxxxxx: _out=147;              //23713536-23713663
                32'b00000001011010011101011110xxxxxx: _out=147;              //23713664-23713727
                32'b00000001011010011101011111000xxx: _out=147;              //23713728-23713735
                32'b0000000101101001110101111100100x: _out=147;              //23713736-23713737
                
                32'b0000000101101001110101111100101x: _out=148;              //23713738-23713739
                32'b000000010110100111010111110011xx: _out=148;              //23713740-23713743
                32'b0000000101101001110101111101xxxx: _out=148;              //23713744-23713759
                32'b000000010110100111010111111xxxxx: _out=148;              //23713760-23713791
                32'b000000010110100111011xxxxxxxxxxx: _out=148;              //23713792-23715839
                32'b0000000101101001111xxxxxxxxxxxxx: _out=148;              //23715840-23724031
                32'b000000010110101xxxxxxxxxxxxxxxxx: _out=148;              //23724032-23855103
                32'b00000001011011xxxxxxxxxxxxxxxxxx: _out=148;              //23855104-24117247
                32'b000000010111xxxxxxxxxxxxxxxxxxxx: _out=148;              //24117248-25165823
                32'b000000011000xxxxxxxxxxxxxxxxxxxx: _out=148;              //25165824-26214399
                32'b00000001100100xxxxxxxxxxxxxxxxxx: _out=148;              //26214400-26476543
                32'b0000000110010100xxxxxxxxxxxxxxxx: _out=148;              //26476544-26542079
                32'b00000001100101010xxxxxxxxxxxxxxx: _out=148;              //26542080-26574847
                32'b000000011001010110xxxxxxxxxxxxxx: _out=148;              //26574848-26591231
                32'b0000000110010101110xxxxxxxxxxxxx: _out=148;              //26591232-26599423
                32'b00000001100101011110xxxxxxxxxxxx: _out=148;              //26599424-26603519
                32'b000000011001010111110xxxxxxxxxxx: _out=148;              //26603520-26605567
                32'b0000000110010101111110xxxxxxxxxx: _out=148;              //26605568-26606591
                32'b00000001100101011111110xxxxxxxxx: _out=148;              //26606592-26607103
                32'b0000000110010101111111100xxxxxxx: _out=148;              //26607104-26607231
                32'b0000000110010101111111101000xxxx: _out=148;              //26607232-26607247
                32'b0000000110010101111111101001000x: _out=148;              //26607248-26607249
                32'b00000001100101011111111010010010: _out=148;              //26607250
                
                32'b00000001100101011111111010010011: _out=149;              //26607251
                32'b000000011001010111111110100101xx: _out=149;              //26607252-26607255
                32'b00000001100101011111111010011xxx: _out=149;              //26607256-26607263
                32'b000000011001010111111110101xxxxx: _out=149;              //26607264-26607295
                32'b00000001100101011111111011xxxxxx: _out=149;              //26607296-26607359
                32'b000000011001010111111111xxxxxxxx: _out=149;              //26607360-26607615
                32'b000000011001011xxxxxxxxxxxxxxxxx: _out=149;              //26607616-26738687
                32'b0000000110011xxxxxxxxxxxxxxxxxxx: _out=149;              //26738688-27262975
                32'b00000001101xxxxxxxxxxxxxxxxxxxxx: _out=149;              //27262976-29360127
                32'b00000001110000xxxxxxxxxxxxxxxxxx: _out=149;              //29360128-29622271
                32'b000000011100010xxxxxxxxxxxxxxxxx: _out=149;              //29622272-29753343
                32'b0000000111000110xxxxxxxxxxxxxxxx: _out=149;              //29753344-29818879
                32'b00000001110001110xxxxxxxxxxxxxxx: _out=149;              //29818880-29851647
                32'b000000011100011110000xxxxxxxxxxx: _out=149;              //29851648-29853695
                32'b0000000111000111100010000xxxxxxx: _out=149;              //29853696-29853823
                32'b0000000111000111100010001000000x: _out=149;              //29853824-29853825
                32'b00000001110001111000100010000010: _out=149;              //29853826
                
                32'b00000001110001111000100010000011: _out=150;              //29853827
                32'b000000011100011110001000100001xx: _out=150;              //29853828-29853831
                32'b00000001110001111000100010001xxx: _out=150;              //29853832-29853839
                32'b0000000111000111100010001001xxxx: _out=150;              //29853840-29853855
                32'b000000011100011110001000101xxxxx: _out=150;              //29853856-29853887
                32'b00000001110001111000100011xxxxxx: _out=150;              //29853888-29853951
                32'b000000011100011110001001xxxxxxxx: _out=150;              //29853952-29854207
                32'b00000001110001111000101xxxxxxxxx: _out=150;              //29854208-29854719
                32'b0000000111000111100011xxxxxxxxxx: _out=150;              //29854720-29855743
                32'b00000001110001111001xxxxxxxxxxxx: _out=150;              //29855744-29859839
                32'b0000000111000111101xxxxxxxxxxxxx: _out=150;              //29859840-29868031
                32'b000000011100011111xxxxxxxxxxxxxx: _out=150;              //29868032-29884415
                32'b0000000111001xxxxxxxxxxxxxxxxxxx: _out=150;              //29884416-30408703
                32'b000000011101xxxxxxxxxxxxxxxxxxxx: _out=150;              //30408704-31457279
                32'b000000011110xxxxxxxxxxxxxxxxxxxx: _out=150;              //31457280-32505855
                32'b0000000111110xxxxxxxxxxxxxxxxxxx: _out=150;              //32505856-33030143
                32'b00000001111110xxxxxxxxxxxxxxxxxx: _out=150;              //33030144-33292287
                32'b000000011111110xxxxxxxxxxxxxxxxx: _out=150;              //33292288-33423359
                32'b0000000111111110xxxxxxxxxxxxxxxx: _out=150;              //33423360-33488895
                32'b00000001111111110000xxxxxxxxxxxx: _out=150;              //33488896-33492991
                32'b000000011111111100010xxxxxxxxxxx: _out=150;              //33492992-33495039
                32'b0000000111111111000110xxxxxxxxxx: _out=150;              //33495040-33496063
                32'b000000011111111100011100xxxxxxxx: _out=150;              //33496064-33496319
                32'b0000000111111111000111010xxxxxxx: _out=150;              //33496320-33496447
                32'b00000001111111110001110110xxxxxx: _out=150;              //33496448-33496511
                32'b000000011111111100011101110xxxxx: _out=150;              //33496512-33496543
                
                32'b000000011111111100011101111xxxxx: _out=151;              //33496544-33496575
                32'b00000001111111110001111xxxxxxxxx: _out=151;              //33496576-33497087
                32'b0000000111111111001xxxxxxxxxxxxx: _out=151;              //33497088-33505279
                32'b000000011111111101xxxxxxxxxxxxxx: _out=151;              //33505280-33521663
                32'b00000001111111111xxxxxxxxxxxxxxx: _out=151;              //33521664-33554431
                32'b00000010000xxxxxxxxxxxxxxxxxxxxx: _out=151;              //33554432-35651583
                32'b000000100010xxxxxxxxxxxxxxxxxxxx: _out=151;              //35651584-36700159
                32'b0000001000110xxxxxxxxxxxxxxxxxxx: _out=151;              //36700160-37224447
                32'b00000010001110xxxxxxxxxxxxxxxxxx: _out=151;              //37224448-37486591
                32'b0000001000111100xxxxxxxxxxxxxxxx: _out=151;              //37486592-37552127
                32'b000000100011110100xxxxxxxxxxxxxx: _out=151;              //37552128-37568511
                32'b0000001000111101010xxxxxxxxxxxxx: _out=151;              //37568512-37576703
                32'b00000010001111010110xxxxxxxxxxxx: _out=151;              //37576704-37580799
                32'b000000100011110101110xxxxxxxxxxx: _out=151;              //37580800-37582847
                32'b00000010001111010111100xxxxxxxxx: _out=151;              //37582848-37583359
                32'b000000100011110101111010xxxxxxxx: _out=151;              //37583360-37583615
                32'b00000010001111010111101100xxxxxx: _out=151;              //37583616-37583679
                32'b000000100011110101111011010xxxxx: _out=151;              //37583680-37583711
                32'b0000001000111101011110110110xxxx: _out=151;              //37583712-37583727
                32'b00000010001111010111101101110xxx: _out=151;              //37583728-37583735
                32'b000000100011110101111011011110xx: _out=151;              //37583736-37583739
                32'b00000010001111010111101101111100: _out=151;              //37583740
                
                32'b00000010001111010111101101111101: _out=152;              //37583741
                32'b0000001000111101011110110111111x: _out=152;              //37583742-37583743
                32'b0000001000111101011110111xxxxxxx: _out=152;              //37583744-37583871
                32'b0000001000111101011111xxxxxxxxxx: _out=152;              //37583872-37584895
                32'b00000010001111011xxxxxxxxxxxxxxx: _out=152;              //37584896-37617663
                32'b000000100011111xxxxxxxxxxxxxxxxx: _out=152;              //37617664-37748735
                32'b0000001001xxxxxxxxxxxxxxxxxxxxxx: _out=152;              //37748736-41943039
                32'b000000101000000xxxxxxxxxxxxxxxxx: _out=152;              //41943040-42074111
                32'b0000001010000010xxxxxxxxxxxxxxxx: _out=152;              //42074112-42139647
                32'b000000101000001100xxxxxxxxxxxxxx: _out=152;              //42139648-42156031
                32'b0000001010000011010xxxxxxxxxxxxx: _out=152;              //42156032-42164223
                32'b00000010100000110110xxxxxxxxxxxx: _out=152;              //42164224-42168319
                32'b0000001010000011011100xxxxxxxxxx: _out=152;              //42168320-42169343
                32'b000000101000001101110100xxxxxxxx: _out=152;              //42169344-42169599
                32'b000000101000001101110101000xxxxx: _out=152;              //42169600-42169631
                32'b0000001010000011011101010010xxxx: _out=152;              //42169632-42169647
                32'b0000001010000011011101010011000x: _out=152;              //42169648-42169649
                32'b00000010100000110111010100110010: _out=152;              //42169650
                
                32'b00000010100000110111010100110011: _out=153;              //42169651
                32'b000000101000001101110101001101xx: _out=153;              //42169652-42169655
                32'b00000010100000110111010100111xxx: _out=153;              //42169656-42169663
                32'b00000010100000110111010101xxxxxx: _out=153;              //42169664-42169727
                32'b0000001010000011011101011xxxxxxx: _out=153;              //42169728-42169855
                32'b00000010100000110111011xxxxxxxxx: _out=153;              //42169856-42170367
                32'b000000101000001101111xxxxxxxxxxx: _out=153;              //42170368-42172415
                32'b00000010100000111xxxxxxxxxxxxxxx: _out=153;              //42172416-42205183
                32'b00000010100001xxxxxxxxxxxxxxxxxx: _out=153;              //42205184-42467327
                32'b0000001010001xxxxxxxxxxxxxxxxxxx: _out=153;              //42467328-42991615
                32'b000000101001xxxxxxxxxxxxxxxxxxxx: _out=153;              //42991616-44040191
                32'b00000010101xxxxxxxxxxxxxxxxxxxxx: _out=153;              //44040192-46137343
                32'b000000101100xxxxxxxxxxxxxxxxxxxx: _out=153;              //46137344-47185919
                32'b0000001011010000xxxxxxxxxxxxxxxx: _out=153;              //47185920-47251455
                32'b00000010110100010xxxxxxxxxxxxxxx: _out=153;              //47251456-47284223
                32'b000000101101000110xxxxxxxxxxxxxx: _out=153;              //47284224-47300607
                32'b0000001011010001110xxxxxxxxxxxxx: _out=153;              //47300608-47308799
                32'b00000010110100011110xxxxxxxxxxxx: _out=153;              //47308800-47312895
                32'b000000101101000111110xxxxxxxxxxx: _out=153;              //47312896-47314943
                32'b0000001011010001111110000xxxxxxx: _out=153;              //47314944-47315071
                32'b000000101101000111111000100xxxxx: _out=153;              //47315072-47315103
                32'b0000001011010001111110001010xxxx: _out=153;              //47315104-47315119
                32'b000000101101000111111000101100xx: _out=153;              //47315120-47315123
                32'b0000001011010001111110001011010x: _out=153;              //47315124-47315125
                
                32'b0000001011010001111110001011011x: _out=154;              //47315126-47315127
                32'b00000010110100011111100010111xxx: _out=154;              //47315128-47315135
                32'b00000010110100011111100011xxxxxx: _out=154;              //47315136-47315199
                32'b000000101101000111111001xxxxxxxx: _out=154;              //47315200-47315455
                32'b00000010110100011111101xxxxxxxxx: _out=154;              //47315456-47315967
                32'b0000001011010001111111xxxxxxxxxx: _out=154;              //47315968-47316991
                32'b000000101101001xxxxxxxxxxxxxxxxx: _out=154;              //47316992-47448063
                32'b00000010110101xxxxxxxxxxxxxxxxxx: _out=154;              //47448064-47710207
                32'b0000001011011xxxxxxxxxxxxxxxxxxx: _out=154;              //47710208-48234495
                32'b00000010111xxxxxxxxxxxxxxxxxxxxx: _out=154;              //48234496-50331647
                32'b00000011000xxxxxxxxxxxxxxxxxxxxx: _out=154;              //50331648-52428799
                32'b0000001100100xxxxxxxxxxxxxxxxxxx: _out=154;              //52428800-52953087
                32'b000000110010100xxxxxxxxxxxxxxxxx: _out=154;              //52953088-53084159
                32'b00000011001010100000xxxxxxxxxxxx: _out=154;              //53084160-53088255
                32'b0000001100101010000100000xxxxxxx: _out=154;              //53088256-53088383
                32'b000000110010101000010000100xxxxx: _out=154;              //53088384-53088415
                32'b0000001100101010000100001010xxxx: _out=154;              //53088416-53088431
                32'b00000011001010100001000010110xxx: _out=154;              //53088432-53088439
                32'b000000110010101000010000101110xx: _out=154;              //53088440-53088443
                32'b00000011001010100001000010111100: _out=154;              //53088444
                
                32'b00000011001010100001000010111101: _out=155;              //53088445
                32'b0000001100101010000100001011111x: _out=155;              //53088446-53088447
                32'b00000011001010100001000011xxxxxx: _out=155;              //53088448-53088511
                32'b000000110010101000010001xxxxxxxx: _out=155;              //53088512-53088767
                32'b00000011001010100001001xxxxxxxxx: _out=155;              //53088768-53089279
                32'b0000001100101010000101xxxxxxxxxx: _out=155;              //53089280-53090303
                32'b000000110010101000011xxxxxxxxxxx: _out=155;              //53090304-53092351
                32'b0000001100101010001xxxxxxxxxxxxx: _out=155;              //53092352-53100543
                32'b000000110010101001xxxxxxxxxxxxxx: _out=155;              //53100544-53116927
                32'b00000011001010101xxxxxxxxxxxxxxx: _out=155;              //53116928-53149695
                32'b0000001100101011xxxxxxxxxxxxxxxx: _out=155;              //53149696-53215231
                32'b00000011001011xxxxxxxxxxxxxxxxxx: _out=155;              //53215232-53477375
                32'b000000110011xxxxxxxxxxxxxxxxxxxx: _out=155;              //53477376-54525951
                32'b0000001101xxxxxxxxxxxxxxxxxxxxxx: _out=155;              //54525952-58720255
                32'b0000001110000xxxxxxxxxxxxxxxxxxx: _out=155;              //58720256-59244543
                32'b00000011100010xxxxxxxxxxxxxxxxxx: _out=155;              //59244544-59506687
                32'b00000011100011000xxxxxxxxxxxxxxx: _out=155;              //59506688-59539455
                32'b000000111000110010xxxxxxxxxxxxxx: _out=155;              //59539456-59555839
                32'b0000001110001100110xxxxxxxxxxxxx: _out=155;              //59555840-59564031
                32'b000000111000110011100xxxxxxxxxxx: _out=155;              //59564032-59566079
                32'b0000001110001100111010000xxxxxxx: _out=155;              //59566080-59566207
                32'b000000111000110011101000100000xx: _out=155;              //59566208-59566211
                32'b0000001110001100111010001000010x: _out=155;              //59566212-59566213
                32'b00000011100011001110100010000110: _out=155;              //59566214
                
                32'b00000011100011001110100010000111: _out=156;              //59566215
                32'b00000011100011001110100010001xxx: _out=156;              //59566216-59566223
                32'b0000001110001100111010001001xxxx: _out=156;              //59566224-59566239
                32'b000000111000110011101000101xxxxx: _out=156;              //59566240-59566271
                32'b00000011100011001110100011xxxxxx: _out=156;              //59566272-59566335
                32'b000000111000110011101001xxxxxxxx: _out=156;              //59566336-59566591
                32'b00000011100011001110101xxxxxxxxx: _out=156;              //59566592-59567103
                32'b0000001110001100111011xxxxxxxxxx: _out=156;              //59567104-59568127
                32'b00000011100011001111xxxxxxxxxxxx: _out=156;              //59568128-59572223
                32'b0000001110001101xxxxxxxxxxxxxxxx: _out=156;              //59572224-59637759
                32'b000000111000111xxxxxxxxxxxxxxxxx: _out=156;              //59637760-59768831
                32'b000000111001xxxxxxxxxxxxxxxxxxxx: _out=156;              //59768832-60817407
                32'b00000011101xxxxxxxxxxxxxxxxxxxxx: _out=156;              //60817408-62914559
                32'b00000011110xxxxxxxxxxxxxxxxxxxxx: _out=156;              //62914560-65011711
                32'b000000111110xxxxxxxxxxxxxxxxxxxx: _out=156;              //65011712-66060287
                32'b0000001111110xxxxxxxxxxxxxxxxxxx: _out=156;              //66060288-66584575
                32'b000000111111100xxxxxxxxxxxxxxxxx: _out=156;              //66584576-66715647
                32'b0000001111111010xxxxxxxxxxxxxxxx: _out=156;              //66715648-66781183
                32'b00000011111110110xxxxxxxxxxxxxxx: _out=156;              //66781184-66813951
                32'b000000111111101110xxxxxxxxxxxxxx: _out=156;              //66813952-66830335
                32'b000000111111101111000xxxxxxxxxxx: _out=156;              //66830336-66832383
                32'b0000001111111011110010xxxxxxxxxx: _out=156;              //66832384-66833407
                32'b00000011111110111100110xxxxxxxxx: _out=156;              //66833408-66833919
                32'b000000111111101111001110xxxxxxxx: _out=156;              //66833920-66834175
                32'b0000001111111011110011110xxxxxxx: _out=156;              //66834176-66834303
                32'b00000011111110111100111110xxxxxx: _out=156;              //66834304-66834367
                32'b0000001111111011110011111100xxxx: _out=156;              //66834368-66834383
                32'b00000011111110111100111111010xxx: _out=156;              //66834384-66834391
                
                32'b00000011111110111100111111011xxx: _out=157;              //66834392-66834399
                32'b000000111111101111001111111xxxxx: _out=157;              //66834400-66834431
                32'b00000011111110111101xxxxxxxxxxxx: _out=157;              //66834432-66838527
                32'b0000001111111011111xxxxxxxxxxxxx: _out=157;              //66838528-66846719
                32'b00000011111111xxxxxxxxxxxxxxxxxx: _out=157;              //66846720-67108863
                32'b0000010000xxxxxxxxxxxxxxxxxxxxxx: _out=157;              //67108864-71303167
                32'b00000100010xxxxxxxxxxxxxxxxxxxxx: _out=157;              //71303168-73400319
                32'b000001000110xxxxxxxxxxxxxxxxxxxx: _out=157;              //73400320-74448895
                32'b0000010001110xxxxxxxxxxxxxxxxxxx: _out=157;              //74448896-74973183
                32'b0000010001111000000xxxxxxxxxxxxx: _out=157;              //74973184-74981375
                32'b00000100011110000010xxxxxxxxxxxx: _out=157;              //74981376-74985471
                32'b000001000111100000110xxxxxxxxxxx: _out=157;              //74985472-74987519
                32'b0000010001111000001110xxxxxxxxxx: _out=157;              //74987520-74988543
                32'b00000100011110000011110xxxxxxxxx: _out=157;              //74988544-74989055
                32'b000001000111100000111110xxxxxxxx: _out=157;              //74989056-74989311
                32'b00000100011110000011111100xxxxxx: _out=157;              //74989312-74989375
                32'b000001000111100000111111010xxxxx: _out=157;              //74989376-74989407
                32'b00000100011110000011111101100xxx: _out=157;              //74989408-74989415
                32'b000001000111100000111111011010xx: _out=157;              //74989416-74989419
                32'b00000100011110000011111101101100: _out=157;              //74989420
                
                32'b00000100011110000011111101101101: _out=158;              //74989421
                32'b0000010001111000001111110110111x: _out=158;              //74989422-74989423
                32'b0000010001111000001111110111xxxx: _out=158;              //74989424-74989439
                32'b0000010001111000001111111xxxxxxx: _out=158;              //74989440-74989567
                32'b000001000111100001xxxxxxxxxxxxxx: _out=158;              //74989568-75005951
                32'b00000100011110001xxxxxxxxxxxxxxx: _out=158;              //75005952-75038719
                32'b0000010001111001xxxxxxxxxxxxxxxx: _out=158;              //75038720-75104255
                32'b000001000111101xxxxxxxxxxxxxxxxx: _out=158;              //75104256-75235327
                32'b00000100011111xxxxxxxxxxxxxxxxxx: _out=158;              //75235328-75497471
                32'b000001001xxxxxxxxxxxxxxxxxxxxxxx: _out=158;              //75497472-83886079
                32'b000001010000000xxxxxxxxxxxxxxxxx: _out=158;              //83886080-84017151
                32'b0000010100000010xxxxxxxxxxxxxxxx: _out=158;              //84017152-84082687
                32'b00000101000000110xxxxxxxxxxxxxxx: _out=158;              //84082688-84115455
                32'b000001010000001110xxxxxxxxxxxxxx: _out=158;              //84115456-84131839
                32'b00000101000000111100xxxxxxxxxxxx: _out=158;              //84131840-84135935
                32'b000001010000001111010xxxxxxxxxxx: _out=158;              //84135936-84137983
                32'b0000010100000011110110xxxxxxxxxx: _out=158;              //84137984-84139007
                32'b000001010000001111011100xxxxxxxx: _out=158;              //84139008-84139263
                32'b0000010100000011110111010xxxxxxx: _out=158;              //84139264-84139391
                32'b00000101000000111101110110xxxxxx: _out=158;              //84139392-84139455
                32'b000001010000001111011101110xxxxx: _out=158;              //84139456-84139487
                32'b0000010100000011110111011110xxxx: _out=158;              //84139488-84139503
                32'b00000101000000111101110111110xxx: _out=158;              //84139504-84139511
                32'b0000010100000011110111011111100x: _out=158;              //84139512-84139513
                32'b00000101000000111101110111111010: _out=158;              //84139514
                
                32'b00000101000000111101110111111011: _out=159;              //84139515
                32'b000001010000001111011101111111xx: _out=159;              //84139516-84139519
                32'b00000101000000111101111xxxxxxxxx: _out=159;              //84139520-84140031
                32'b0000010100000011111xxxxxxxxxxxxx: _out=159;              //84140032-84148223
                32'b00000101000001xxxxxxxxxxxxxxxxxx: _out=159;              //84148224-84410367
                32'b0000010100001xxxxxxxxxxxxxxxxxxx: _out=159;              //84410368-84934655
                32'b000001010001xxxxxxxxxxxxxxxxxxxx: _out=159;              //84934656-85983231
                32'b00000101001xxxxxxxxxxxxxxxxxxxxx: _out=159;              //85983232-88080383
                32'b0000010101xxxxxxxxxxxxxxxxxxxxxx: _out=159;              //88080384-92274687
                32'b00000101100xxxxxxxxxxxxxxxxxxxxx: _out=159;              //92274688-94371839
                32'b00000101101000000xxxxxxxxxxxxxxx: _out=159;              //94371840-94404607
                32'b0000010110100000100000xxxxxxxxxx: _out=159;              //94404608-94405631
                32'b000001011010000010000100xxxxxxxx: _out=159;              //94405632-94405887
                32'b0000010110100000100001010xxxxxxx: _out=159;              //94405888-94406015
                32'b00000101101000001000010110xxxxxx: _out=159;              //94406016-94406079
                32'b00000101101000001000010111000xxx: _out=159;              //94406080-94406087
                
                32'b00000101101000001000010111001xxx: _out=160;              //94406088-94406095
                32'b0000010110100000100001011101xxxx: _out=160;              //94406096-94406111
                32'b000001011010000010000101111xxxxx: _out=160;              //94406112-94406143
                32'b00000101101000001000011xxxxxxxxx: _out=160;              //94406144-94406655
                32'b000001011010000010001xxxxxxxxxxx: _out=160;              //94406656-94408703
                32'b00000101101000001001xxxxxxxxxxxx: _out=160;              //94408704-94412799
                32'b0000010110100000101xxxxxxxxxxxxx: _out=160;              //94412800-94420991
                32'b000001011010000011xxxxxxxxxxxxxx: _out=160;              //94420992-94437375
                32'b0000010110100001xxxxxxxxxxxxxxxx: _out=160;              //94437376-94502911
                32'b000001011010001xxxxxxxxxxxxxxxxx: _out=160;              //94502912-94633983
                32'b00000101101001xxxxxxxxxxxxxxxxxx: _out=160;              //94633984-94896127
                32'b0000010110101xxxxxxxxxxxxxxxxxxx: _out=160;              //94896128-95420415
                32'b000001011011xxxxxxxxxxxxxxxxxxxx: _out=160;              //95420416-96468991
                32'b0000010111xxxxxxxxxxxxxxxxxxxxxx: _out=160;              //96468992-100663295
                32'b0000011000xxxxxxxxxxxxxxxxxxxxxx: _out=160;              //100663296-104857599
                32'b000001100100xxxxxxxxxxxxxxxxxxxx: _out=160;              //104857600-105906175
                32'b000001100101000000xxxxxxxxxxxxxx: _out=160;              //105906176-105922559
                32'b000001100101000001000xxxxxxxxxxx: _out=160;              //105922560-105924607
                32'b00000110010100000100100xxxxxxxxx: _out=160;              //105924608-105925119
                32'b0000011001010000010010100xxxxxxx: _out=160;              //105925120-105925247
                32'b00000110010100000100101010xxxxxx: _out=160;              //105925248-105925311
                32'b000001100101000001001010110xxxxx: _out=160;              //105925312-105925343
                32'b0000011001010000010010101110xxxx: _out=160;              //105925344-105925359
                32'b00000110010100000100101011110xxx: _out=160;              //105925360-105925367
                32'b000001100101000001001010111110xx: _out=160;              //105925368-105925371
                32'b00000110010100000100101011111100: _out=160;              //105925372
                
                32'b00000110010100000100101011111101: _out=161;              //105925373
                32'b0000011001010000010010101111111x: _out=161;              //105925374-105925375
                32'b000001100101000001001011xxxxxxxx: _out=161;              //105925376-105925631
                32'b0000011001010000010011xxxxxxxxxx: _out=161;              //105925632-105926655
                32'b00000110010100000101xxxxxxxxxxxx: _out=161;              //105926656-105930751
                32'b0000011001010000011xxxxxxxxxxxxx: _out=161;              //105930752-105938943
                32'b00000110010100001xxxxxxxxxxxxxxx: _out=161;              //105938944-105971711
                32'b0000011001010001xxxxxxxxxxxxxxxx: _out=161;              //105971712-106037247
                32'b000001100101001xxxxxxxxxxxxxxxxx: _out=161;              //106037248-106168319
                32'b00000110010101xxxxxxxxxxxxxxxxxx: _out=161;              //106168320-106430463
                32'b0000011001011xxxxxxxxxxxxxxxxxxx: _out=161;              //106430464-106954751
                32'b00000110011xxxxxxxxxxxxxxxxxxxxx: _out=161;              //106954752-109051903
                32'b000001101xxxxxxxxxxxxxxxxxxxxxxx: _out=161;              //109051904-117440511
                32'b000001110000xxxxxxxxxxxxxxxxxxxx: _out=161;              //117440512-118489087
                32'b00000111000100xxxxxxxxxxxxxxxxxx: _out=161;              //118489088-118751231
                32'b0000011100010100xxxxxxxxxxxxxxxx: _out=161;              //118751232-118816767
                32'b00000111000101010xxxxxxxxxxxxxxx: _out=161;              //118816768-118849535
                32'b00000111000101011000000xxxxxxxxx: _out=161;              //118849536-118850047
                32'b0000011100010101100000100xxxxxxx: _out=161;              //118850048-118850175
                32'b000001110001010110000010100xxxxx: _out=161;              //118850176-118850207
                32'b00000111000101011000001010100xxx: _out=161;              //118850208-118850215
                32'b000001110001010110000010101010xx: _out=161;              //118850216-118850219
                32'b0000011100010101100000101010110x: _out=161;              //118850220-118850221
                32'b00000111000101011000001010101110: _out=161;              //118850222
                
                32'b00000111000101011000001010101111: _out=162;              //118850223
                32'b0000011100010101100000101011xxxx: _out=162;              //118850224-118850239
                32'b00000111000101011000001011xxxxxx: _out=162;              //118850240-118850303
                32'b000001110001010110000011xxxxxxxx: _out=162;              //118850304-118850559
                32'b0000011100010101100001xxxxxxxxxx: _out=162;              //118850560-118851583
                32'b000001110001010110001xxxxxxxxxxx: _out=162;              //118851584-118853631
                32'b00000111000101011001xxxxxxxxxxxx: _out=162;              //118853632-118857727
                32'b0000011100010101101xxxxxxxxxxxxx: _out=162;              //118857728-118865919
                32'b000001110001010111xxxxxxxxxxxxxx: _out=162;              //118865920-118882303
                32'b000001110001011xxxxxxxxxxxxxxxxx: _out=162;              //118882304-119013375
                32'b0000011100011xxxxxxxxxxxxxxxxxxx: _out=162;              //119013376-119537663
                32'b00000111001xxxxxxxxxxxxxxxxxxxxx: _out=162;              //119537664-121634815
                32'b0000011101xxxxxxxxxxxxxxxxxxxxxx: _out=162;              //121634816-125829119
                32'b0000011110xxxxxxxxxxxxxxxxxxxxxx: _out=162;              //125829120-130023423
                32'b00000111110xxxxxxxxxxxxxxxxxxxxx: _out=162;              //130023424-132120575
                32'b000001111110xxxxxxxxxxxxxxxxxxxx: _out=162;              //132120576-133169151
                32'b000001111111000xxxxxxxxxxxxxxxxx: _out=162;              //133169152-133300223
                32'b00000111111100100xxxxxxxxxxxxxxx: _out=162;              //133300224-133332991
                32'b000001111111001010xxxxxxxxxxxxxx: _out=162;              //133332992-133349375
                32'b000001111111001011000xxxxxxxxxxx: _out=162;              //133349376-133351423
                32'b00000111111100101100100xxxxxxxxx: _out=162;              //133351424-133351935
                32'b0000011111110010110010100xxxxxxx: _out=162;              //133351936-133352063
                32'b00000111111100101100101010xxxxxx: _out=162;              //133352064-133352127
                32'b0000011111110010110010101100xxxx: _out=162;              //133352128-133352143
                
                32'b0000011111110010110010101101xxxx: _out=163;              //133352144-133352159
                32'b000001111111001011001010111xxxxx: _out=163;              //133352160-133352191
                32'b000001111111001011001011xxxxxxxx: _out=163;              //133352192-133352447
                32'b0000011111110010110011xxxxxxxxxx: _out=163;              //133352448-133353471
                32'b00000111111100101101xxxxxxxxxxxx: _out=163;              //133353472-133357567
                32'b0000011111110010111xxxxxxxxxxxxx: _out=163;              //133357568-133365759
                32'b0000011111110011xxxxxxxxxxxxxxxx: _out=163;              //133365760-133431295
                32'b00000111111101xxxxxxxxxxxxxxxxxx: _out=163;              //133431296-133693439
                32'b0000011111111xxxxxxxxxxxxxxxxxxx: _out=163;              //133693440-134217727
                32'b000010000xxxxxxxxxxxxxxxxxxxxxxx: _out=163;              //134217728-142606335
                32'b0000100010xxxxxxxxxxxxxxxxxxxxxx: _out=163;              //142606336-146800639
                32'b00001000110xxxxxxxxxxxxxxxxxxxxx: _out=163;              //146800640-148897791
                32'b0000100011100xxxxxxxxxxxxxxxxxxx: _out=163;              //148897792-149422079
                32'b000010001110100xxxxxxxxxxxxxxxxx: _out=163;              //149422080-149553151
                32'b0000100011101010xxxxxxxxxxxxxxxx: _out=163;              //149553152-149618687
                32'b00001000111010110000xxxxxxxxxxxx: _out=163;              //149618688-149622783
                32'b00001000111010110001000xxxxxxxxx: _out=163;              //149622784-149623295
                32'b000010001110101100010010xxxxxxxx: _out=163;              //149623296-149623551
                32'b00001000111010110001001100000xxx: _out=163;              //149623552-149623559
                32'b000010001110101100010011000010xx: _out=163;              //149623560-149623563
                32'b0000100011101011000100110000110x: _out=163;              //149623564-149623565
                
                32'b0000100011101011000100110000111x: _out=164;              //149623566-149623567
                32'b0000100011101011000100110001xxxx: _out=164;              //149623568-149623583
                32'b000010001110101100010011001xxxxx: _out=164;              //149623584-149623615
                32'b00001000111010110001001101xxxxxx: _out=164;              //149623616-149623679
                32'b0000100011101011000100111xxxxxxx: _out=164;              //149623680-149623807
                32'b0000100011101011000101xxxxxxxxxx: _out=164;              //149623808-149624831
                32'b000010001110101100011xxxxxxxxxxx: _out=164;              //149624832-149626879
                32'b0000100011101011001xxxxxxxxxxxxx: _out=164;              //149626880-149635071
                32'b000010001110101101xxxxxxxxxxxxxx: _out=164;              //149635072-149651455
                32'b00001000111010111xxxxxxxxxxxxxxx: _out=164;              //149651456-149684223
                32'b00001000111011xxxxxxxxxxxxxxxxxx: _out=164;              //149684224-149946367
                32'b000010001111xxxxxxxxxxxxxxxxxxxx: _out=164;              //149946368-150994943
                32'b00001001xxxxxxxxxxxxxxxxxxxxxxxx: _out=164;              //150994944-167772159
                32'b0000101000000000xxxxxxxxxxxxxxxx: _out=164;              //167772160-167837695
                32'b00001010000000010xxxxxxxxxxxxxxx: _out=164;              //167837696-167870463
                32'b0000101000000001100xxxxxxxxxxxxx: _out=164;              //167870464-167878655
                32'b0000101000000001101000xxxxxxxxxx: _out=164;              //167878656-167879679
                32'b00001010000000011010010xxxxxxxxx: _out=164;              //167879680-167880191
                32'b0000101000000001101001100xxxxxxx: _out=164;              //167880192-167880319
                32'b00001010000000011010011010xxxxxx: _out=164;              //167880320-167880383
                32'b0000101000000001101001101100xxxx: _out=164;              //167880384-167880399
                32'b0000101000000001101001101101000x: _out=164;              //167880400-167880401
                
                32'b0000101000000001101001101101001x: _out=165;              //167880402-167880403
                32'b000010100000000110100110110101xx: _out=165;              //167880404-167880407
                32'b00001010000000011010011011011xxx: _out=165;              //167880408-167880415
                32'b000010100000000110100110111xxxxx: _out=165;              //167880416-167880447
                32'b000010100000000110100111xxxxxxxx: _out=165;              //167880448-167880703
                32'b000010100000000110101xxxxxxxxxxx: _out=165;              //167880704-167882751
                32'b00001010000000011011xxxxxxxxxxxx: _out=165;              //167882752-167886847
                32'b000010100000000111xxxxxxxxxxxxxx: _out=165;              //167886848-167903231
                32'b000010100000001xxxxxxxxxxxxxxxxx: _out=165;              //167903232-168034303
                32'b00001010000001xxxxxxxxxxxxxxxxxx: _out=165;              //168034304-168296447
                32'b0000101000001xxxxxxxxxxxxxxxxxxx: _out=165;              //168296448-168820735
                32'b000010100001xxxxxxxxxxxxxxxxxxxx: _out=165;              //168820736-169869311
                32'b00001010001xxxxxxxxxxxxxxxxxxxxx: _out=165;              //169869312-171966463
                32'b0000101001xxxxxxxxxxxxxxxxxxxxxx: _out=165;              //171966464-176160767
                32'b000010101xxxxxxxxxxxxxxxxxxxxxxx: _out=165;              //176160768-184549375
                32'b00001011000xxxxxxxxxxxxxxxxxxxxx: _out=165;              //184549376-186646527
                32'b000010110010xxxxxxxxxxxxxxxxxxxx: _out=165;              //186646528-187695103
                32'b0000101100110xxxxxxxxxxxxxxxxxxx: _out=165;              //187695104-188219391
                32'b000010110011100xxxxxxxxxxxxxxxxx: _out=165;              //188219392-188350463
                32'b0000101100111010000xxxxxxxxxxxxx: _out=165;              //188350464-188358655
                32'b00001011001110100010xxxxxxxxxxxx: _out=165;              //188358656-188362751
                32'b000010110011101000110xxxxxxxxxxx: _out=165;              //188362752-188364799
                32'b00001011001110100011100000xxxxxx: _out=165;              //188364800-188364863
                32'b000010110011101000111000010xxxxx: _out=165;              //188364864-188364895
                32'b00001011001110100011100001100xxx: _out=165;              //188364896-188364903
                32'b000010110011101000111000011010xx: _out=165;              //188364904-188364907
                32'b00001011001110100011100001101100: _out=165;              //188364908
                
                32'b00001011001110100011100001101101: _out=166;              //188364909
                32'b0000101100111010001110000110111x: _out=166;              //188364910-188364911
                32'b0000101100111010001110000111xxxx: _out=166;              //188364912-188364927
                32'b0000101100111010001110001xxxxxxx: _out=166;              //188364928-188365055
                32'b000010110011101000111001xxxxxxxx: _out=166;              //188365056-188365311
                32'b00001011001110100011101xxxxxxxxx: _out=166;              //188365312-188365823
                32'b0000101100111010001111xxxxxxxxxx: _out=166;              //188365824-188366847
                32'b000010110011101001xxxxxxxxxxxxxx: _out=166;              //188366848-188383231
                32'b00001011001110101xxxxxxxxxxxxxxx: _out=166;              //188383232-188415999
                32'b0000101100111011xxxxxxxxxxxxxxxx: _out=166;              //188416000-188481535
                32'b00001011001111xxxxxxxxxxxxxxxxxx: _out=166;              //188481536-188743679
                32'b0000101101xxxxxxxxxxxxxxxxxxxxxx: _out=166;              //188743680-192937983
                32'b000010111xxxxxxxxxxxxxxxxxxxxxxx: _out=166;              //192937984-201326591
                32'b000011000xxxxxxxxxxxxxxxxxxxxxxx: _out=166;              //201326592-209715199
                32'b000011001000xxxxxxxxxxxxxxxxxxxx: _out=166;              //209715200-210763775
                32'b0000110010010xxxxxxxxxxxxxxxxxxx: _out=166;              //210763776-211288063
                32'b00001100100110000xxxxxxxxxxxxxxx: _out=166;              //211288064-211320831
                32'b000011001001100010xxxxxxxxxxxxxx: _out=166;              //211320832-211337215
                32'b0000110010011000110xxxxxxxxxxxxx: _out=166;              //211337216-211345407
                32'b000011001001100011100xxxxxxxxxxx: _out=166;              //211345408-211347455
                32'b0000110010011000111010xxxxxxxxxx: _out=166;              //211347456-211348479
                32'b000011001001100011101100xxxxxxxx: _out=166;              //211348480-211348735
                32'b0000110010011000111011010xxxxxxx: _out=166;              //211348736-211348863
                32'b000011001001100011101101100xxxxx: _out=166;              //211348864-211348895
                32'b00001100100110001110110110100xxx: _out=166;              //211348896-211348903
                
                32'b00001100100110001110110110101xxx: _out=167;              //211348904-211348911
                32'b0000110010011000111011011011xxxx: _out=167;              //211348912-211348927
                32'b00001100100110001110110111xxxxxx: _out=167;              //211348928-211348991
                32'b00001100100110001110111xxxxxxxxx: _out=167;              //211348992-211349503
                32'b00001100100110001111xxxxxxxxxxxx: _out=167;              //211349504-211353599
                32'b0000110010011001xxxxxxxxxxxxxxxx: _out=167;              //211353600-211419135
                32'b000011001001101xxxxxxxxxxxxxxxxx: _out=167;              //211419136-211550207
                32'b00001100100111xxxxxxxxxxxxxxxxxx: _out=167;              //211550208-211812351
                32'b00001100101xxxxxxxxxxxxxxxxxxxxx: _out=167;              //211812352-213909503
                32'b0000110011xxxxxxxxxxxxxxxxxxxxxx: _out=167;              //213909504-218103807
                32'b00001101xxxxxxxxxxxxxxxxxxxxxxxx: _out=167;              //218103808-234881023
                32'b00001110000xxxxxxxxxxxxxxxxxxxxx: _out=167;              //234881024-236978175
                32'b000011100010000xxxxxxxxxxxxxxxxx: _out=167;              //236978176-237109247
                32'b000011100010001000xxxxxxxxxxxxxx: _out=167;              //237109248-237125631
                32'b0000111000100010010xxxxxxxxxxxxx: _out=167;              //237125632-237133823
                32'b000011100010001001100xxxxxxxxxxx: _out=167;              //237133824-237135871
                32'b0000111000100010011010xxxxxxxxxx: _out=167;              //237135872-237136895
                32'b000011100010001001101100xxxxxxxx: _out=167;              //237136896-237137151
                32'b0000111000100010011011010xxxxxxx: _out=167;              //237137152-237137279
                32'b00001110001000100110110110xxxxxx: _out=167;              //237137280-237137343
                32'b0000111000100010011011011100xxxx: _out=167;              //237137344-237137359
                32'b00001110001000100110110111010xxx: _out=167;              //237137360-237137367
                32'b0000111000100010011011011101100x: _out=167;              //237137368-237137369
                32'b00001110001000100110110111011010: _out=167;              //237137370
                
                32'b00001110001000100110110111011011: _out=168;              //237137371
                32'b000011100010001001101101110111xx: _out=168;              //237137372-237137375
                32'b000011100010001001101101111xxxxx: _out=168;              //237137376-237137407
                32'b00001110001000100110111xxxxxxxxx: _out=168;              //237137408-237137919
                32'b00001110001000100111xxxxxxxxxxxx: _out=168;              //237137920-237142015
                32'b00001110001000101xxxxxxxxxxxxxxx: _out=168;              //237142016-237174783
                32'b0000111000100011xxxxxxxxxxxxxxxx: _out=168;              //237174784-237240319
                32'b00001110001001xxxxxxxxxxxxxxxxxx: _out=168;              //237240320-237502463
                32'b0000111000101xxxxxxxxxxxxxxxxxxx: _out=168;              //237502464-238026751
                32'b000011100011xxxxxxxxxxxxxxxxxxxx: _out=168;              //238026752-239075327
                32'b0000111001xxxxxxxxxxxxxxxxxxxxxx: _out=168;              //239075328-243269631
                32'b000011101xxxxxxxxxxxxxxxxxxxxxxx: _out=168;              //243269632-251658239
                32'b000011110xxxxxxxxxxxxxxxxxxxxxxx: _out=168;              //251658240-260046847
                32'b0000111110xxxxxxxxxxxxxxxxxxxxxx: _out=168;              //260046848-264241151
                32'b000011111100xxxxxxxxxxxxxxxxxxxx: _out=168;              //264241152-265289727
                32'b0000111111010xxxxxxxxxxxxxxxxxxx: _out=168;              //265289728-265814015
                32'b000011111101100xxxxxxxxxxxxxxxxx: _out=168;              //265814016-265945087
                32'b0000111111011010xxxxxxxxxxxxxxxx: _out=168;              //265945088-266010623
                32'b00001111110110110xxxxxxxxxxxxxxx: _out=168;              //266010624-266043391
                32'b000011111101101110xxxxxxxxxxxxxx: _out=168;              //266043392-266059775
                32'b0000111111011011110xxxxxxxxxxxxx: _out=168;              //266059776-266067967
                32'b00001111110110111110xxxxxxxxxxxx: _out=168;              //266067968-266072063
                32'b000011111101101111110000xxxxxxxx: _out=168;              //266072064-266072319
                32'b0000111111011011111100010xxxxxxx: _out=168;              //266072320-266072447
                32'b000011111101101111110001100xxxxx: _out=168;              //266072448-266072479
                32'b0000111111011011111100011010xxxx: _out=168;              //266072480-266072495
                32'b00001111110110111111000110110xxx: _out=168;              //266072496-266072503
                32'b0000111111011011111100011011100x: _out=168;              //266072504-266072505
                
                32'b0000111111011011111100011011101x: _out=169;              //266072506-266072507
                32'b000011111101101111110001101111xx: _out=169;              //266072508-266072511
                32'b00001111110110111111000111xxxxxx: _out=169;              //266072512-266072575
                32'b00001111110110111111001xxxxxxxxx: _out=169;              //266072576-266073087
                32'b0000111111011011111101xxxxxxxxxx: _out=169;              //266073088-266074111
                32'b000011111101101111111xxxxxxxxxxx: _out=169;              //266074112-266076159
                32'b00001111110111xxxxxxxxxxxxxxxxxx: _out=169;              //266076160-266338303
                32'b00001111111xxxxxxxxxxxxxxxxxxxxx: _out=169;              //266338304-268435455
                32'b00010000xxxxxxxxxxxxxxxxxxxxxxxx: _out=169;              //268435456-285212671
                32'b000100010xxxxxxxxxxxxxxxxxxxxxxx: _out=169;              //285212672-293601279
                32'b0001000110xxxxxxxxxxxxxxxxxxxxxx: _out=169;              //293601280-297795583
                32'b0001000111000xxxxxxxxxxxxxxxxxxx: _out=169;              //297795584-298319871
                32'b000100011100100xxxxxxxxxxxxxxxxx: _out=169;              //298319872-298450943
                32'b0001000111001010xxxxxxxxxxxxxxxx: _out=169;              //298450944-298516479
                32'b000100011100101100xxxxxxxxxxxxxx: _out=169;              //298516480-298532863
                32'b00010001110010110100xxxxxxxxxxxx: _out=169;              //298532864-298536959
                32'b0001000111001011010100xxxxxxxxxx: _out=169;              //298536960-298537983
                32'b000100011100101101010100xxxxxxxx: _out=169;              //298537984-298538239
                32'b0001000111001011010101010000xxxx: _out=169;              //298538240-298538255
                32'b000100011100101101010101000100xx: _out=169;              //298538256-298538259
                32'b0001000111001011010101010001010x: _out=169;              //298538260-298538261
                
                32'b0001000111001011010101010001011x: _out=170;              //298538262-298538263
                32'b00010001110010110101010100011xxx: _out=170;              //298538264-298538271
                32'b000100011100101101010101001xxxxx: _out=170;              //298538272-298538303
                32'b00010001110010110101010101xxxxxx: _out=170;              //298538304-298538367
                32'b0001000111001011010101011xxxxxxx: _out=170;              //298538368-298538495
                32'b00010001110010110101011xxxxxxxxx: _out=170;              //298538496-298539007
                32'b000100011100101101011xxxxxxxxxxx: _out=170;              //298539008-298541055
                32'b0001000111001011011xxxxxxxxxxxxx: _out=170;              //298541056-298549247
                32'b00010001110010111xxxxxxxxxxxxxxx: _out=170;              //298549248-298582015
                32'b00010001110011xxxxxxxxxxxxxxxxxx: _out=170;              //298582016-298844159
                32'b000100011101xxxxxxxxxxxxxxxxxxxx: _out=170;              //298844160-299892735
                32'b00010001111xxxxxxxxxxxxxxxxxxxxx: _out=170;              //299892736-301989887
                32'b00010010xxxxxxxxxxxxxxxxxxxxxxxx: _out=170;              //301989888-318767103
                32'b000100110xxxxxxxxxxxxxxxxxxxxxxx: _out=170;              //318767104-327155711
                32'b0001001110xxxxxxxxxxxxxxxxxxxxxx: _out=170;              //327155712-331350015
                32'b00010011110xxxxxxxxxxxxxxxxxxxxx: _out=170;              //331350016-333447167
                32'b000100111110xxxxxxxxxxxxxxxxxxxx: _out=170;              //333447168-334495743
                32'b00010011111100xxxxxxxxxxxxxxxxxx: _out=170;              //334495744-334757887
                32'b000100111111010xxxxxxxxxxxxxxxxx: _out=170;              //334757888-334888959
                32'b0001001111110110xxxxxxxxxxxxxxxx: _out=170;              //334888960-334954495
                32'b0001001111110111000xxxxxxxxxxxxx: _out=170;              //334954496-334962687
                32'b000100111111011100100xxxxxxxxxxx: _out=170;              //334962688-334964735
                32'b00010011111101110010100xxxxxxxxx: _out=170;              //334964736-334965247
                32'b0001001111110111001010100xxxxxxx: _out=170;              //334965248-334965375
                32'b00010011111101110010101010xxxxxx: _out=170;              //334965376-334965439

                32'b00010011111101110010101011xxxxxx: _out=171;              //334965440-334965503
                32'b000100111111011100101011xxxxxxxx: _out=171;              //334965504-334965759
                32'b0001001111110111001011xxxxxxxxxx: _out=171;              //334965760-334966783
                32'b00010011111101110011xxxxxxxxxxxx: _out=171;              //334966784-334970879
                32'b000100111111011101xxxxxxxxxxxxxx: _out=171;              //334970880-334987263
                32'b00010011111101111xxxxxxxxxxxxxxx: _out=171;              //334987264-335020031
                32'b0001001111111xxxxxxxxxxxxxxxxxxx: _out=171;              //335020032-335544319
                32'b0001010xxxxxxxxxxxxxxxxxxxxxxxxx: _out=171;              //335544320-369098751
                32'b0001011000xxxxxxxxxxxxxxxxxxxxxx: _out=171;              //369098752-373293055
                32'b00010110010xxxxxxxxxxxxxxxxxxxxx: _out=171;              //373293056-375390207
                32'b00010110011000xxxxxxxxxxxxxxxxxx: _out=171;              //375390208-375652351
                32'b000101100110010xxxxxxxxxxxxxxxxx: _out=171;              //375652352-375783423
                32'b00010110011001100xxxxxxxxxxxxxxx: _out=171;              //375783424-375816191
                32'b000101100110011010xxxxxxxxxxxxxx: _out=171;              //375816192-375832575
                32'b00010110011001101100xxxxxxxxxxxx: _out=171;              //375832576-375836671
                32'b00010110011001101101000xxxxxxxxx: _out=171;              //375836672-375837183
                32'b0001011001100110110100100xxxxxxx: _out=171;              //375837184-375837311
                32'b00010110011001101101001010xxxxxx: _out=171;              //375837312-375837375
                32'b0001011001100110110100101100xxxx: _out=171;              //375837376-375837391
                32'b00010110011001101101001011010xxx: _out=171;              //375837392-375837399
                32'b000101100110011011010010110110xx: _out=171;              //375837400-375837403
                32'b00010110011001101101001011011100: _out=171;              //375837404
                
                32'b00010110011001101101001011011101: _out=172;              //375837405
                32'b0001011001100110110100101101111x: _out=172;              //375837406-375837407
                32'b000101100110011011010010111xxxxx: _out=172;              //375837408-375837439
                32'b000101100110011011010011xxxxxxxx: _out=172;              //375837440-375837695
                32'b0001011001100110110101xxxxxxxxxx: _out=172;              //375837696-375838719
                32'b000101100110011011011xxxxxxxxxxx: _out=172;              //375838720-375840767
                32'b0001011001100110111xxxxxxxxxxxxx: _out=172;              //375840768-375848959
                32'b0001011001100111xxxxxxxxxxxxxxxx: _out=172;              //375848960-375914495
                32'b0001011001101xxxxxxxxxxxxxxxxxxx: _out=172;              //375914496-376438783
                32'b000101100111xxxxxxxxxxxxxxxxxxxx: _out=172;              //376438784-377487359
                32'b000101101xxxxxxxxxxxxxxxxxxxxxxx: _out=172;              //377487360-385875967
                32'b00010111xxxxxxxxxxxxxxxxxxxxxxxx: _out=172;              //385875968-402653183
                32'b00011000xxxxxxxxxxxxxxxxxxxxxxxx: _out=172;              //402653184-419430399
                32'b00011001000xxxxxxxxxxxxxxxxxxxxx: _out=172;              //419430400-421527551
                32'b000110010010000xxxxxxxxxxxxxxxxx: _out=172;              //421527552-421658623
                32'b00011001001000100xxxxxxxxxxxxxxx: _out=172;              //421658624-421691391
                32'b00011001001000101000xxxxxxxxxxxx: _out=172;              //421691392-421695487
                32'b00011001001000101001000xxxxxxxxx: _out=172;              //421695488-421695999
                32'b000110010010001010010010xxxxxxxx: _out=172;              //421696000-421696255
                32'b0001100100100010100100110xxxxxxx: _out=172;              //421696256-421696383
                32'b00011001001000101001001110xxxxxx: _out=172;              //421696384-421696447
                32'b000110010010001010010011110xxxxx: _out=172;              //421696448-421696479
                32'b0001100100100010100100111110xxxx: _out=172;              //421696480-421696495
                32'b00011001001000101001001111110xxx: _out=172;              //421696496-421696503
                
                32'b00011001001000101001001111111xxx: _out=173;              //421696504-421696511
                32'b0001100100100010100101xxxxxxxxxx: _out=173;              //421696512-421697535
                32'b000110010010001010011xxxxxxxxxxx: _out=173;              //421697536-421699583
                32'b0001100100100010101xxxxxxxxxxxxx: _out=173;              //421699584-421707775
                32'b000110010010001011xxxxxxxxxxxxxx: _out=173;              //421707776-421724159
                32'b0001100100100011xxxxxxxxxxxxxxxx: _out=173;              //421724160-421789695
                32'b00011001001001xxxxxxxxxxxxxxxxxx: _out=173;              //421789696-422051839
                32'b0001100100101xxxxxxxxxxxxxxxxxxx: _out=173;              //422051840-422576127
                32'b000110010011xxxxxxxxxxxxxxxxxxxx: _out=173;              //422576128-423624703
                32'b0001100101xxxxxxxxxxxxxxxxxxxxxx: _out=173;              //423624704-427819007
                32'b000110011xxxxxxxxxxxxxxxxxxxxxxx: _out=173;              //427819008-436207615
                32'b0001101xxxxxxxxxxxxxxxxxxxxxxxxx: _out=173;              //436207616-469762047
                32'b00011100000xxxxxxxxxxxxxxxxxxxxx: _out=173;              //469762048-471859199
                32'b000111000010xxxxxxxxxxxxxxxxxxxx: _out=173;              //471859200-472907775
                32'b000111000011000xxxxxxxxxxxxxxxxx: _out=173;              //472907776-473038847
                32'b0001110000110010xxxxxxxxxxxxxxxx: _out=173;              //473038848-473104383
                32'b00011100001100110xxxxxxxxxxxxxxx: _out=173;              //473104384-473137151
                32'b0001110000110011100xxxxxxxxxxxxx: _out=173;              //473137152-473145343
                32'b00011100001100111010xxxxxxxxxxxx: _out=173;              //473145344-473149439
                32'b0001110000110011101100xxxxxxxxxx: _out=173;              //473149440-473150463
                32'b00011100001100111011010xxxxxxxxx: _out=173;              //473150464-473150975
                32'b000111000011001110110110xxxxxxxx: _out=173;              //473150976-473151231
                32'b0001110000110011101101110000xxxx: _out=173;              //473151232-473151247
                32'b00011100001100111011011100010xxx: _out=173;              //473151248-473151255
                32'b0001110000110011101101110001100x: _out=173;              //473151256-473151257
                32'b00011100001100111011011100011010: _out=173;              //473151258
                
                32'b00011100001100111011011100011011: _out=174;              //473151259
                32'b000111000011001110110111000111xx: _out=174;              //473151260-473151263
                32'b000111000011001110110111001xxxxx: _out=174;              //473151264-473151295
                32'b00011100001100111011011101xxxxxx: _out=174;              //473151296-473151359
                32'b0001110000110011101101111xxxxxxx: _out=174;              //473151360-473151487
                32'b000111000011001110111xxxxxxxxxxx: _out=174;              //473151488-473153535
                32'b000111000011001111xxxxxxxxxxxxxx: _out=174;              //473153536-473169919
                32'b00011100001101xxxxxxxxxxxxxxxxxx: _out=174;              //473169920-473432063
                32'b0001110000111xxxxxxxxxxxxxxxxxxx: _out=174;              //473432064-473956351
                32'b0001110001xxxxxxxxxxxxxxxxxxxxxx: _out=174;              //473956352-478150655
                32'b000111001xxxxxxxxxxxxxxxxxxxxxxx: _out=174;              //478150656-486539263
                32'b00011101xxxxxxxxxxxxxxxxxxxxxxxx: _out=174;              //486539264-503316479
                32'b00011110xxxxxxxxxxxxxxxxxxxxxxxx: _out=174;              //503316480-520093695
                32'b000111110xxxxxxxxxxxxxxxxxxxxxxx: _out=174;              //520093696-528482303
                32'b00011111100xxxxxxxxxxxxxxxxxxxxx: _out=174;              //528482304-530579455
                32'b00011111101000xxxxxxxxxxxxxxxxxx: _out=174;              //530579456-530841599
                32'b00011111101001000xxxxxxxxxxxxxxx: _out=174;              //530841600-530874367
                32'b0001111110100100100xxxxxxxxxxxxx: _out=174;              //530874368-530882559
                32'b0001111110100100101000xxxxxxxxxx: _out=174;              //530882560-530883583
                32'b00011111101001001010010xxxxxxxxx: _out=174;              //530883584-530884095
                32'b000111111010010010100110xxxxxxxx: _out=174;              //530884096-530884351
                32'b00011111101001001010011100xxxxxx: _out=174;              //530884352-530884415
                32'b0001111110100100101001110100xxxx: _out=174;              //530884416-530884431
                32'b00011111101001001010011101010xxx: _out=174;              //530884432-530884439
                32'b000111111010010010100111010110xx: _out=174;              //530884440-530884443
                32'b00011111101001001010011101011100: _out=174;              //530884444
                
                32'b00011111101001001010011101011101: _out=175;              //530884445
                32'b0001111110100100101001110101111x: _out=175;              //530884446-530884447
                32'b000111111010010010100111011xxxxx: _out=175;              //530884448-530884479
                32'b0001111110100100101001111xxxxxxx: _out=175;              //530884480-530884607
                32'b000111111010010010101xxxxxxxxxxx: _out=175;              //530884608-530886655
                32'b00011111101001001011xxxxxxxxxxxx: _out=175;              //530886656-530890751
                32'b000111111010010011xxxxxxxxxxxxxx: _out=175;              //530890752-530907135
                32'b0001111110100101xxxxxxxxxxxxxxxx: _out=175;              //530907136-530972671
                32'b000111111010011xxxxxxxxxxxxxxxxx: _out=175;              //530972672-531103743
                32'b0001111110101xxxxxxxxxxxxxxxxxxx: _out=175;              //531103744-531628031
                32'b000111111011xxxxxxxxxxxxxxxxxxxx: _out=175;              //531628032-532676607
                32'b0001111111xxxxxxxxxxxxxxxxxxxxxx: _out=175;              //532676608-536870911
                32'b0010000xxxxxxxxxxxxxxxxxxxxxxxxx: _out=175;              //536870912-570425343
                32'b00100010xxxxxxxxxxxxxxxxxxxxxxxx: _out=175;              //570425344-587202559
                32'b001000110xxxxxxxxxxxxxxxxxxxxxxx: _out=175;              //587202560-595591167
                32'b0010001110000000xxxxxxxxxxxxxxxx: _out=175;              //595591168-595656703
                32'b00100011100000010000xxxxxxxxxxxx: _out=175;              //595656704-595660799
                32'b0010001110000001000100xxxxxxxxxx: _out=175;              //595660800-595661823
                32'b001000111000000100010100xxxxxxxx: _out=175;              //595661824-595662079
                32'b00100011100000010001010100xxxxxx: _out=175;              //595662080-595662143
                
                32'b00100011100000010001010101xxxxxx: _out=176;              //595662144-595662207
                32'b0010001110000001000101011xxxxxxx: _out=176;              //595662208-595662335
                32'b00100011100000010001011xxxxxxxxx: _out=176;              //595662336-595662847
                32'b001000111000000100011xxxxxxxxxxx: _out=176;              //595662848-595664895
                32'b0010001110000001001xxxxxxxxxxxxx: _out=176;              //595664896-595673087
                32'b001000111000000101xxxxxxxxxxxxxx: _out=176;              //595673088-595689471
                32'b00100011100000011xxxxxxxxxxxxxxx: _out=176;              //595689472-595722239
                32'b001000111000001xxxxxxxxxxxxxxxxx: _out=176;              //595722240-595853311
                32'b00100011100001xxxxxxxxxxxxxxxxxx: _out=176;              //595853312-596115455
                32'b0010001110001xxxxxxxxxxxxxxxxxxx: _out=176;              //596115456-596639743
                32'b001000111001xxxxxxxxxxxxxxxxxxxx: _out=176;              //596639744-597688319
                32'b00100011101xxxxxxxxxxxxxxxxxxxxx: _out=176;              //597688320-599785471
                32'b0010001111xxxxxxxxxxxxxxxxxxxxxx: _out=176;              //599785472-603979775
                32'b0010010xxxxxxxxxxxxxxxxxxxxxxxxx: _out=176;              //603979776-637534207
                32'b00100110xxxxxxxxxxxxxxxxxxxxxxxx: _out=176;              //637534208-654311423
                32'b001001110xxxxxxxxxxxxxxxxxxxxxxx: _out=176;              //654311424-662700031
                32'b0010011110xxxxxxxxxxxxxxxxxxxxxx: _out=176;              //662700032-666894335
                32'b001001111100xxxxxxxxxxxxxxxxxxxx: _out=176;              //666894336-667942911
                32'b00100111110100xxxxxxxxxxxxxxxxxx: _out=176;              //667942912-668205055
                32'b001001111101010xxxxxxxxxxxxxxxxx: _out=176;              //668205056-668336127
                32'b00100111110101100000xxxxxxxxxxxx: _out=176;              //668336128-668340223
                32'b001001111101011000010xxxxxxxxxxx: _out=176;              //668340224-668342271
                32'b0010011111010110000110xxxxxxxxxx: _out=176;              //668342272-668343295
                32'b00100111110101100001110xxxxxxxxx: _out=176;              //668343296-668343807
                32'b00100111110101100001111000xxxxxx: _out=176;              //668343808-668343871
                32'b001001111101011000011110010xxxxx: _out=176;              //668343872-668343903
                32'b00100111110101100001111001100xxx: _out=176;              //668343904-668343911
                32'b001001111101011000011110011010xx: _out=176;              //668343912-668343915
                32'b0010011111010110000111100110110x: _out=176;              //668343916-668343917
                
                32'b0010011111010110000111100110111x: _out=177;              //668343918-668343919
                32'b0010011111010110000111100111xxxx: _out=177;              //668343920-668343935
                32'b0010011111010110000111101xxxxxxx: _out=177;              //668343936-668344063
                32'b001001111101011000011111xxxxxxxx: _out=177;              //668344064-668344319
                32'b0010011111010110001xxxxxxxxxxxxx: _out=177;              //668344320-668352511
                32'b001001111101011001xxxxxxxxxxxxxx: _out=177;              //668352512-668368895
                32'b00100111110101101xxxxxxxxxxxxxxx: _out=177;              //668368896-668401663
                32'b0010011111010111xxxxxxxxxxxxxxxx: _out=177;              //668401664-668467199
                32'b0010011111011xxxxxxxxxxxxxxxxxxx: _out=177;              //668467200-668991487
                32'b00100111111xxxxxxxxxxxxxxxxxxxxx: _out=177;              //668991488-671088639
                32'b001010xxxxxxxxxxxxxxxxxxxxxxxxxx: _out=177;              //671088640-738197503
                32'b001011000xxxxxxxxxxxxxxxxxxxxxxx: _out=177;              //738197504-746586111
                32'b00101100100xxxxxxxxxxxxxxxxxxxxx: _out=177;              //746586112-748683263
                32'b001011001010xxxxxxxxxxxxxxxxxxxx: _out=177;              //748683264-749731839
                32'b001011001011000xxxxxxxxxxxxxxxxx: _out=177;              //749731840-749862911
                32'b001011001011001000xxxxxxxxxxxxxx: _out=177;              //749862912-749879295
                32'b0010110010110010010xxxxxxxxxxxxx: _out=177;              //749879296-749887487
                32'b00101100101100100110xxxxxxxxxxxx: _out=177;              //749887488-749891583
                32'b001011001011001001110xxxxxxxxxxx: _out=177;              //749891584-749893631
                32'b00101100101100100111100xxxxxxxxx: _out=177;              //749893632-749894143
                32'b00101100101100100111101000xxxxxx: _out=177;              //749894144-749894207
                32'b0010110010110010011110100100000x: _out=177;              //749894208-749894209
                
                32'b0010110010110010011110100100001x: _out=178;              //749894210-749894211
                32'b001011001011001001111010010001xx: _out=178;              //749894212-749894215
                32'b00101100101100100111101001001xxx: _out=178;              //749894216-749894223
                32'b0010110010110010011110100101xxxx: _out=178;              //749894224-749894239
                32'b001011001011001001111010011xxxxx: _out=178;              //749894240-749894271
                32'b0010110010110010011110101xxxxxxx: _out=178;              //749894272-749894399
                32'b001011001011001001111011xxxxxxxx: _out=178;              //749894400-749894655
                32'b0010110010110010011111xxxxxxxxxx: _out=178;              //749894656-749895679
                32'b00101100101100101xxxxxxxxxxxxxxx: _out=178;              //749895680-749928447
                32'b0010110010110011xxxxxxxxxxxxxxxx: _out=178;              //749928448-749993983
                32'b00101100101101xxxxxxxxxxxxxxxxxx: _out=178;              //749993984-750256127
                32'b0010110010111xxxxxxxxxxxxxxxxxxx: _out=178;              //750256128-750780415
                32'b0010110011xxxxxxxxxxxxxxxxxxxxxx: _out=178;              //750780416-754974719
                32'b00101101xxxxxxxxxxxxxxxxxxxxxxxx: _out=178;              //754974720-771751935
                32'b0010111xxxxxxxxxxxxxxxxxxxxxxxxx: _out=178;              //771751936-805306367
                32'b0011000xxxxxxxxxxxxxxxxxxxxxxxxx: _out=178;              //805306368-838860799
                32'b00110010000xxxxxxxxxxxxxxxxxxxxx: _out=178;              //838860800-840957951
                32'b00110010001000xxxxxxxxxxxxxxxxxx: _out=178;              //840957952-841220095
                32'b001100100010010xxxxxxxxxxxxxxxxx: _out=178;              //841220096-841351167
                32'b00110010001001100xxxxxxxxxxxxxxx: _out=178;              //841351168-841383935
                32'b0011001000100110100xxxxxxxxxxxxx: _out=178;              //841383936-841392127
                32'b001100100010011010100xxxxxxxxxxx: _out=178;              //841392128-841394175
                32'b00110010001001101010100xxxxxxxxx: _out=178;              //841394176-841394687
                32'b001100100010011010101010xxxxxxxx: _out=178;              //841394688-841394943
                32'b0011001000100110101010110xxxxxxx: _out=178;              //841394944-841395071
                32'b00110010001001101010101110xxxxxx: _out=178;              //841395072-841395135
                32'b001100100010011010101011110000xx: _out=178;              //841395136-841395139
                32'b0011001000100110101010111100010x: _out=178;              //841395140-841395141
                
                32'b0011001000100110101010111100011x: _out=179;              //841395142-841395143
                32'b00110010001001101010101111001xxx: _out=179;              //841395144-841395151
                32'b0011001000100110101010111101xxxx: _out=179;              //841395152-841395167
                32'b001100100010011010101011111xxxxx: _out=179;              //841395168-841395199
                32'b0011001000100110101011xxxxxxxxxx: _out=179;              //841395200-841396223
                32'b00110010001001101011xxxxxxxxxxxx: _out=179;              //841396224-841400319
                32'b001100100010011011xxxxxxxxxxxxxx: _out=179;              //841400320-841416703
                32'b0011001000100111xxxxxxxxxxxxxxxx: _out=179;              //841416704-841482239
                32'b0011001000101xxxxxxxxxxxxxxxxxxx: _out=179;              //841482240-842006527
                32'b001100100011xxxxxxxxxxxxxxxxxxxx: _out=179;              //842006528-843055103
                32'b0011001001xxxxxxxxxxxxxxxxxxxxxx: _out=179;              //843055104-847249407
                32'b001100101xxxxxxxxxxxxxxxxxxxxxxx: _out=179;              //847249408-855638015
                32'b00110011xxxxxxxxxxxxxxxxxxxxxxxx: _out=179;              //855638016-872415231
                32'b001101xxxxxxxxxxxxxxxxxxxxxxxxxx: _out=179;              //872415232-939524095
                32'b0011100000xxxxxxxxxxxxxxxxxxxxxx: _out=179;              //939524096-943718399
                32'b00111000010000xxxxxxxxxxxxxxxxxx: _out=179;              //943718400-943980543
                32'b0011100001000100xxxxxxxxxxxxxxxx: _out=179;              //943980544-944046079
                32'b0011100001000101000xxxxxxxxxxxxx: _out=179;              //944046080-944054271
                32'b00111000010001010010xxxxxxxxxxxx: _out=179;              //944054272-944058367
                32'b001110000100010100110xxxxxxxxxxx: _out=179;              //944058368-944060415
                32'b001110000100010100111000xxxxxxxx: _out=179;              //944060416-944060671
                32'b0011100001000101001110010xxxxxxx: _out=179;              //944060672-944060799
                32'b00111000010001010011100110xxxxxx: _out=179;              //944060800-944060863
                32'b00111000010001010011100111000xxx: _out=179;              //944060864-944060871
                32'b001110000100010100111001110010xx: _out=179;              //944060872-944060875
                32'b00111000010001010011100111001100: _out=179;              //944060876
                
                32'b00111000010001010011100111001101: _out=180;              //944060877
                32'b0011100001000101001110011100111x: _out=180;              //944060878-944060879
                32'b0011100001000101001110011101xxxx: _out=180;              //944060880-944060895
                32'b001110000100010100111001111xxxxx: _out=180;              //944060896-944060927
                32'b00111000010001010011101xxxxxxxxx: _out=180;              //944060928-944061439
                32'b0011100001000101001111xxxxxxxxxx: _out=180;              //944061440-944062463
                32'b001110000100010101xxxxxxxxxxxxxx: _out=180;              //944062464-944078847
                32'b00111000010001011xxxxxxxxxxxxxxx: _out=180;              //944078848-944111615
                32'b001110000100011xxxxxxxxxxxxxxxxx: _out=180;              //944111616-944242687
                32'b0011100001001xxxxxxxxxxxxxxxxxxx: _out=180;              //944242688-944766975
                32'b001110000101xxxxxxxxxxxxxxxxxxxx: _out=180;              //944766976-945815551
                32'b00111000011xxxxxxxxxxxxxxxxxxxxx: _out=180;              //945815552-947912703
                32'b001110001xxxxxxxxxxxxxxxxxxxxxxx: _out=180;              //947912704-956301311
                32'b00111001xxxxxxxxxxxxxxxxxxxxxxxx: _out=180;              //956301312-973078527
                32'b0011101xxxxxxxxxxxxxxxxxxxxxxxxx: _out=180;              //973078528-1006632959
                32'b0011110xxxxxxxxxxxxxxxxxxxxxxxxx: _out=180;              //1006632960-1040187391
                32'b00111110xxxxxxxxxxxxxxxxxxxxxxxx: _out=180;              //1040187392-1056964607
                32'b00111111000xxxxxxxxxxxxxxxxxxxxx: _out=180;              //1056964608-1059061759
                32'b001111110010000xxxxxxxxxxxxxxxxx: _out=180;              //1059061760-1059192831
                32'b00111111001000100xxxxxxxxxxxxxxx: _out=180;              //1059192832-1059225599
                32'b001111110010001010xxxxxxxxxxxxxx: _out=180;              //1059225600-1059241983
                32'b0011111100100010110xxxxxxxxxxxxx: _out=180;              //1059241984-1059250175
                32'b001111110010001011100xxxxxxxxxxx: _out=180;              //1059250176-1059252223
                32'b0011111100100010111010xxxxxxxxxx: _out=180;              //1059252224-1059253247
                32'b001111110010001011101100xxxxxxxx: _out=180;              //1059253248-1059253503
                32'b0011111100100010111011010xxxxxxx: _out=180;              //1059253504-1059253631
                32'b00111111001000101110110110xxxxxx: _out=180;              //1059253632-1059253695
                32'b0011111100100010111011011100xxxx: _out=180;              //1059253696-1059253711
                32'b00111111001000101110110111010xxx: _out=180;              //1059253712-1059253719
                32'b001111110010001011101101110110xx: _out=180;              //1059253720-1059253723
                32'b0011111100100010111011011101110x: _out=180;              //1059253724-1059253725
                
                32'b0011111100100010111011011101111x: _out=181;              //1059253726-1059253727
                32'b001111110010001011101101111xxxxx: _out=181;              //1059253728-1059253759
                32'b00111111001000101110111xxxxxxxxx: _out=181;              //1059253760-1059254271
                32'b00111111001000101111xxxxxxxxxxxx: _out=181;              //1059254272-1059258367
                32'b0011111100100011xxxxxxxxxxxxxxxx: _out=181;              //1059258368-1059323903
                32'b00111111001001xxxxxxxxxxxxxxxxxx: _out=181;              //1059323904-1059586047
                32'b0011111100101xxxxxxxxxxxxxxxxxxx: _out=181;              //1059586048-1060110335
                32'b001111110011xxxxxxxxxxxxxxxxxxxx: _out=181;              //1060110336-1061158911
                32'b0011111101xxxxxxxxxxxxxxxxxxxxxx: _out=181;              //1061158912-1065353215
                32'b001111111xxxxxxxxxxxxxxxxxxxxxxx: _out=181;              //1065353216-1073741823
                32'b010000xxxxxxxxxxxxxxxxxxxxxxxxxx: _out=181;              //1073741824-1140850687
                32'b0100010xxxxxxxxxxxxxxxxxxxxxxxxx: _out=181;              //1140850688-1174405119
                32'b010001100xxxxxxxxxxxxxxxxxxxxxxx: _out=181;              //1174405120-1182793727
                32'b0100011010xxxxxxxxxxxxxxxxxxxxxx: _out=181;              //1182793728-1186988031
                32'b010001101100xxxxxxxxxxxxxxxxxxxx: _out=181;              //1186988032-1188036607
                32'b01000110110100xxxxxxxxxxxxxxxxxx: _out=181;              //1188036608-1188298751
                32'b010001101101010xxxxxxxxxxxxxxxxx: _out=181;              //1188298752-1188429823
                32'b0100011011010110xxxxxxxxxxxxxxxx: _out=181;              //1188429824-1188495359
                32'b01000110110101110000xxxxxxxxxxxx: _out=181;              //1188495360-1188499455
                32'b010001101101011100010xxxxxxxxxxx: _out=181;              //1188499456-1188501503
                32'b01000110110101110001100xxxxxxxxx: _out=181;              //1188501504-1188502015
                32'b0100011011010111000110100xxxxxxx: _out=181;              //1188502016-1188502143
                32'b01000110110101110001101010xxxxxx: _out=181;              //1188502144-1188502207
                32'b0100011011010111000110101100xxxx: _out=181;              //1188502208-1188502223
                32'b010001101101011100011010110100xx: _out=181;              //1188502224-1188502227
                
                32'b010001101101011100011010110101xx: _out=182;              //1188502228-1188502231
                32'b01000110110101110001101011011xxx: _out=182;              //1188502232-1188502239
                32'b010001101101011100011010111xxxxx: _out=182;              //1188502240-1188502271
                32'b010001101101011100011011xxxxxxxx: _out=182;              //1188502272-1188502527
                32'b0100011011010111000111xxxxxxxxxx: _out=182;              //1188502528-1188503551
                32'b0100011011010111001xxxxxxxxxxxxx: _out=182;              //1188503552-1188511743
                32'b010001101101011101xxxxxxxxxxxxxx: _out=182;              //1188511744-1188528127
                32'b01000110110101111xxxxxxxxxxxxxxx: _out=182;              //1188528128-1188560895
                32'b0100011011011xxxxxxxxxxxxxxxxxxx: _out=182;              //1188560896-1189085183
                32'b01000110111xxxxxxxxxxxxxxxxxxxxx: _out=182;              //1189085184-1191182335
                32'b01000111xxxxxxxxxxxxxxxxxxxxxxxx: _out=182;              //1191182336-1207959551
                32'b010010xxxxxxxxxxxxxxxxxxxxxxxxxx: _out=182;              //1207959552-1275068415
                32'b0100110xxxxxxxxxxxxxxxxxxxxxxxxx: _out=182;              //1275068416-1308622847
                32'b01001110xxxxxxxxxxxxxxxxxxxxxxxx: _out=182;              //1308622848-1325400063
                32'b0100111100xxxxxxxxxxxxxxxxxxxxxx: _out=182;              //1325400064-1329594367
                32'b01001111010xxxxxxxxxxxxxxxxxxxxx: _out=182;              //1329594368-1331691519
                32'b010011110110xxxxxxxxxxxxxxxxxxxx: _out=182;              //1331691520-1332740095
                32'b0100111101110xxxxxxxxxxxxxxxxxxx: _out=182;              //1332740096-1333264383
                32'b010011110111100xxxxxxxxxxxxxxxxx: _out=182;              //1333264384-1333395455
                32'b0100111101111010xxxxxxxxxxxxxxxx: _out=182;              //1333395456-1333460991
                32'b01001111011110110xxxxxxxxxxxxxxx: _out=182;              //1333460992-1333493759
                32'b010011110111101110xxxxxxxxxxxxxx: _out=182;              //1333493760-1333510143
                32'b0100111101111011110xxxxxxxxxxxxx: _out=182;              //1333510144-1333518335
                32'b010011110111101111100xxxxxxxxxxx: _out=182;              //1333518336-1333520383
                32'b0100111101111011111010xxxxxxxxxx: _out=182;              //1333520384-1333521407
                32'b0100111101111011111011000000xxxx: _out=182;              //1333521408-1333521423
                32'b01001111011110111110110000010xxx: _out=182;              //1333521424-1333521431
                32'b01001111011110111110110000011000: _out=182;              //1333521432
                
                32'b01001111011110111110110000011001: _out=183;              //1333521433
                32'b0100111101111011111011000001101x: _out=183;              //1333521434-1333521435
                32'b010011110111101111101100000111xx: _out=183;              //1333521436-1333521439
                32'b010011110111101111101100001xxxxx: _out=183;              //1333521440-1333521471
                32'b01001111011110111110110001xxxxxx: _out=183;              //1333521472-1333521535
                32'b0100111101111011111011001xxxxxxx: _out=183;              //1333521536-1333521663
                32'b010011110111101111101101xxxxxxxx: _out=183;              //1333521664-1333521919
                32'b01001111011110111110111xxxxxxxxx: _out=183;              //1333521920-1333522431
                32'b01001111011110111111xxxxxxxxxxxx: _out=183;              //1333522432-1333526527
                32'b01001111011111xxxxxxxxxxxxxxxxxx: _out=183;              //1333526528-1333788671
                32'b010011111xxxxxxxxxxxxxxxxxxxxxxx: _out=183;              //1333788672-1342177279
                32'b01010xxxxxxxxxxxxxxxxxxxxxxxxxxx: _out=183;              //1342177280-1476395007
                32'b01011000xxxxxxxxxxxxxxxxxxxxxxxx: _out=183;              //1476395008-1493172223
                32'b01011001000xxxxxxxxxxxxxxxxxxxxx: _out=183;              //1493172224-1495269375
                32'b0101100100100xxxxxxxxxxxxxxxxxxx: _out=183;              //1495269376-1495793663
                32'b01011001001010xxxxxxxxxxxxxxxxxx: _out=183;              //1495793664-1496055807
                32'b010110010010110xxxxxxxxxxxxxxxxx: _out=183;              //1496055808-1496186879
                32'b01011001001011100xxxxxxxxxxxxxxx: _out=183;              //1496186880-1496219647
                32'b0101100100101110100xxxxxxxxxxxxx: _out=183;              //1496219648-1496227839
                32'b01011001001011101010xxxxxxxxxxxx: _out=183;              //1496227840-1496231935
                32'b010110010010111010110xxxxxxxxxxx: _out=183;              //1496231936-1496233983
                32'b0101100100101110101110xxxxxxxxxx: _out=183;              //1496233984-1496235007
                32'b01011001001011101011110xxxxxxxxx: _out=183;              //1496235008-1496235519
                32'b0101100100101110101111100xxxxxxx: _out=183;              //1496235520-1496235647
                32'b01011001001011101011111010000xxx: _out=183;              //1496235648-1496235655
                32'b01011001001011101011111010001000: _out=183;              //1496235656
                
                32'b01011001001011101011111010001001: _out=184;              //1496235657
                32'b0101100100101110101111101000101x: _out=184;              //1496235658-1496235659
                32'b010110010010111010111110100011xx: _out=184;              //1496235660-1496235663
                32'b0101100100101110101111101001xxxx: _out=184;              //1496235664-1496235679
                32'b010110010010111010111110101xxxxx: _out=184;              //1496235680-1496235711
                32'b01011001001011101011111011xxxxxx: _out=184;              //1496235712-1496235775
                32'b010110010010111010111111xxxxxxxx: _out=184;              //1496235776-1496236031
                32'b010110010010111011xxxxxxxxxxxxxx: _out=184;              //1496236032-1496252415
                32'b0101100100101111xxxxxxxxxxxxxxxx: _out=184;              //1496252416-1496317951
                32'b010110010011xxxxxxxxxxxxxxxxxxxx: _out=184;              //1496317952-1497366527
                32'b0101100101xxxxxxxxxxxxxxxxxxxxxx: _out=184;              //1497366528-1501560831
                32'b010110011xxxxxxxxxxxxxxxxxxxxxxx: _out=184;              //1501560832-1509949439
                32'b0101101xxxxxxxxxxxxxxxxxxxxxxxxx: _out=184;              //1509949440-1543503871
                32'b010111xxxxxxxxxxxxxxxxxxxxxxxxxx: _out=184;              //1543503872-1610612735
                32'b011000xxxxxxxxxxxxxxxxxxxxxxxxxx: _out=184;              //1610612736-1677721599
                32'b011001000000xxxxxxxxxxxxxxxxxxxx: _out=184;              //1677721600-1678770175
                32'b01100100000100000xxxxxxxxxxxxxxx: _out=184;              //1678770176-1678802943
                32'b0110010000010000100000xxxxxxxxxx: _out=184;              //1678802944-1678803967
                32'b011001000001000010000100000xxxxx: _out=184;              //1678803968-1678803999
                32'b0110010000010000100001000010xxxx: _out=184;              //1678804000-1678804015
                32'b0110010000010000100001000011000x: _out=184;              //1678804016-1678804017
                32'b01100100000100001000010000110010: _out=184;              //1678804018
                
                32'b01100100000100001000010000110011: _out=185;              //1678804019
                32'b011001000001000010000100001101xx: _out=185;              //1678804020-1678804023
                32'b01100100000100001000010000111xxx: _out=185;              //1678804024-1678804031
                32'b01100100000100001000010001xxxxxx: _out=185;              //1678804032-1678804095
                32'b0110010000010000100001001xxxxxxx: _out=185;              //1678804096-1678804223
                32'b011001000001000010000101xxxxxxxx: _out=185;              //1678804224-1678804479
                32'b01100100000100001000011xxxxxxxxx: _out=185;              //1678804480-1678804991
                32'b011001000001000010001xxxxxxxxxxx: _out=185;              //1678804992-1678807039
                32'b01100100000100001001xxxxxxxxxxxx: _out=185;              //1678807040-1678811135
                32'b0110010000010000101xxxxxxxxxxxxx: _out=185;              //1678811136-1678819327
                32'b011001000001000011xxxxxxxxxxxxxx: _out=185;              //1678819328-1678835711
                32'b0110010000010001xxxxxxxxxxxxxxxx: _out=185;              //1678835712-1678901247
                32'b011001000001001xxxxxxxxxxxxxxxxx: _out=185;              //1678901248-1679032319
                32'b01100100000101xxxxxxxxxxxxxxxxxx: _out=185;              //1679032320-1679294463
                32'b0110010000011xxxxxxxxxxxxxxxxxxx: _out=185;              //1679294464-1679818751
                32'b01100100001xxxxxxxxxxxxxxxxxxxxx: _out=185;              //1679818752-1681915903
                32'b0110010001xxxxxxxxxxxxxxxxxxxxxx: _out=185;              //1681915904-1686110207
                32'b011001001xxxxxxxxxxxxxxxxxxxxxxx: _out=185;              //1686110208-1694498815
                32'b01100101xxxxxxxxxxxxxxxxxxxxxxxx: _out=185;              //1694498816-1711276031
                32'b0110011xxxxxxxxxxxxxxxxxxxxxxxxx: _out=185;              //1711276032-1744830463
                32'b01101xxxxxxxxxxxxxxxxxxxxxxxxxxx: _out=185;              //1744830464-1879048191
                32'b0111000000xxxxxxxxxxxxxxxxxxxxxx: _out=185;              //1879048192-1883242495
                32'b01110000010000xxxxxxxxxxxxxxxxxx: _out=185;              //1883242496-1883504639
                32'b011100000100010xxxxxxxxxxxxxxxxx: _out=185;              //1883504640-1883635711
                32'b0111000001000110000xxxxxxxxxxxxx: _out=185;              //1883635712-1883643903
                32'b01110000010001100010xxxxxxxxxxxx: _out=185;              //1883643904-1883647999
                32'b0111000001000110001100xxxxxxxxxx: _out=185;              //1883648000-1883649023
                32'b01110000010001100011010000xxxxxx: _out=185;              //1883649024-1883649087
                32'b0111000001000110001101000100000x: _out=185;              //1883649088-1883649089
                
                32'b0111000001000110001101000100001x: _out=186;              //1883649090-1883649091
                32'b011100000100011000110100010001xx: _out=186;              //1883649092-1883649095
                32'b01110000010001100011010001001xxx: _out=186;              //1883649096-1883649103
                32'b0111000001000110001101000101xxxx: _out=186;              //1883649104-1883649119
                32'b011100000100011000110100011xxxxx: _out=186;              //1883649120-1883649151
                32'b0111000001000110001101001xxxxxxx: _out=186;              //1883649152-1883649279
                32'b011100000100011000110101xxxxxxxx: _out=186;              //1883649280-1883649535
                32'b01110000010001100011011xxxxxxxxx: _out=186;              //1883649536-1883650047
                32'b011100000100011000111xxxxxxxxxxx: _out=186;              //1883650048-1883652095
                32'b011100000100011001xxxxxxxxxxxxxx: _out=186;              //1883652096-1883668479
                32'b01110000010001101xxxxxxxxxxxxxxx: _out=186;              //1883668480-1883701247
                32'b0111000001000111xxxxxxxxxxxxxxxx: _out=186;              //1883701248-1883766783
                32'b0111000001001xxxxxxxxxxxxxxxxxxx: _out=186;              //1883766784-1884291071
                32'b011100000101xxxxxxxxxxxxxxxxxxxx: _out=186;              //1884291072-1885339647
                32'b01110000011xxxxxxxxxxxxxxxxxxxxx: _out=186;              //1885339648-1887436799
                32'b011100001xxxxxxxxxxxxxxxxxxxxxxx: _out=186;              //1887436800-1895825407
                32'b01110001xxxxxxxxxxxxxxxxxxxxxxxx: _out=186;              //1895825408-1912602623
                32'b0111001xxxxxxxxxxxxxxxxxxxxxxxxx: _out=186;              //1912602624-1946157055
                32'b011101xxxxxxxxxxxxxxxxxxxxxxxxxx: _out=186;              //1946157056-2013265919
                32'b011110xxxxxxxxxxxxxxxxxxxxxxxxxx: _out=186;              //2013265920-2080374783
                32'b01111100xxxxxxxxxxxxxxxxxxxxxxxx: _out=186;              //2080374784-2097151999
                32'b011111010xxxxxxxxxxxxxxxxxxxxxxx: _out=186;              //2097152000-2105540607
                32'b0111110110xxxxxxxxxxxxxxxxxxxxxx: _out=186;              //2105540608-2109734911
                32'b01111101110xxxxxxxxxxxxxxxxxxxxx: _out=186;              //2109734912-2111832063
                32'b011111011110xxxxxxxxxxxxxxxxxxxx: _out=186;              //2111832064-2112880639
                32'b0111110111110xxxxxxxxxxxxxxxxxxx: _out=186;              //2112880640-2113404927
                32'b0111110111111000xxxxxxxxxxxxxxxx: _out=186;              //2113404928-2113470463
                32'b011111011111100100xxxxxxxxxxxxxx: _out=186;              //2113470464-2113486847
                32'b011111011111100101000xxxxxxxxxxx: _out=186;              //2113486848-2113488895
                32'b0111110111111001010010000xxxxxxx: _out=186;              //2113488896-2113489023
                32'b0111110111111001010010001000xxxx: _out=186;              //2113489024-2113489039
                
                32'b0111110111111001010010001001xxxx: _out=187;              //2113489040-2113489055
                32'b011111011111100101001000101xxxxx: _out=187;              //2113489056-2113489087
                32'b01111101111110010100100011xxxxxx: _out=187;              //2113489088-2113489151
                32'b011111011111100101001001xxxxxxxx: _out=187;              //2113489152-2113489407
                32'b01111101111110010100101xxxxxxxxx: _out=187;              //2113489408-2113489919
                32'b0111110111111001010011xxxxxxxxxx: _out=187;              //2113489920-2113490943
                32'b01111101111110010101xxxxxxxxxxxx: _out=187;              //2113490944-2113495039
                32'b0111110111111001011xxxxxxxxxxxxx: _out=187;              //2113495040-2113503231
                32'b01111101111110011xxxxxxxxxxxxxxx: _out=187;              //2113503232-2113535999
                32'b011111011111101xxxxxxxxxxxxxxxxx: _out=187;              //2113536000-2113667071
                32'b01111101111111xxxxxxxxxxxxxxxxxx: _out=187;              //2113667072-2113929215
                32'b0111111xxxxxxxxxxxxxxxxxxxxxxxxx: _out=187;              //2113929216-2147483647
                32'b10000xxxxxxxxxxxxxxxxxxxxxxxxxxx: _out=187;              //2147483648-2281701375
                32'b100010xxxxxxxxxxxxxxxxxxxxxxxxxx: _out=187;              //2281701376-2348810239
                32'b10001100xxxxxxxxxxxxxxxxxxxxxxxx: _out=187;              //2348810240-2365587455
                32'b1000110100xxxxxxxxxxxxxxxxxxxxxx: _out=187;              //2365587456-2369781759
                32'b100011010100xxxxxxxxxxxxxxxxxxxx: _out=187;              //2369781760-2370830335
                32'b1000110101010xxxxxxxxxxxxxxxxxxx: _out=187;              //2370830336-2371354623
                32'b100011010101100000xxxxxxxxxxxxxx: _out=187;              //2371354624-2371371007
                32'b100011010101100001000xxxxxxxxxxx: _out=187;              //2371371008-2371373055
                32'b10001101010110000100100xxxxxxxxx: _out=187;              //2371373056-2371373567
                32'b1000110101011000010010100xxxxxxx: _out=187;              //2371373568-2371373695
                32'b10001101010110000100101010000xxx: _out=187;              //2371373696-2371373703
                32'b1000110101011000010010101000100x: _out=187;              //2371373704-2371373705
                
                32'b1000110101011000010010101000101x: _out=188;              //2371373706-2371373707
                32'b100011010101100001001010100011xx: _out=188;              //2371373708-2371373711
                32'b1000110101011000010010101001xxxx: _out=188;              //2371373712-2371373727
                32'b100011010101100001001010101xxxxx: _out=188;              //2371373728-2371373759
                32'b10001101010110000100101011xxxxxx: _out=188;              //2371373760-2371373823
                32'b100011010101100001001011xxxxxxxx: _out=188;              //2371373824-2371374079
                32'b1000110101011000010011xxxxxxxxxx: _out=188;              //2371374080-2371375103
                32'b10001101010110000101xxxxxxxxxxxx: _out=188;              //2371375104-2371379199
                32'b1000110101011000011xxxxxxxxxxxxx: _out=188;              //2371379200-2371387391
                32'b10001101010110001xxxxxxxxxxxxxxx: _out=188;              //2371387392-2371420159
                32'b1000110101011001xxxxxxxxxxxxxxxx: _out=188;              //2371420160-2371485695
                32'b100011010101101xxxxxxxxxxxxxxxxx: _out=188;              //2371485696-2371616767
                32'b10001101010111xxxxxxxxxxxxxxxxxx: _out=188;              //2371616768-2371878911
                32'b10001101011xxxxxxxxxxxxxxxxxxxxx: _out=188;              //2371878912-2373976063
                32'b100011011xxxxxxxxxxxxxxxxxxxxxxx: _out=188;              //2373976064-2382364671
                32'b1000111xxxxxxxxxxxxxxxxxxxxxxxxx: _out=188;              //2382364672-2415919103
                32'b10010xxxxxxxxxxxxxxxxxxxxxxxxxxx: _out=188;              //2415919104-2550136831
                32'b100110xxxxxxxxxxxxxxxxxxxxxxxxxx: _out=188;              //2550136832-2617245695
                32'b1001110xxxxxxxxxxxxxxxxxxxxxxxxx: _out=188;              //2617245696-2650800127
                32'b100111100xxxxxxxxxxxxxxxxxxxxxxx: _out=188;              //2650800128-2659188735
                32'b100111101000xxxxxxxxxxxxxxxxxxxx: _out=188;              //2659188736-2660237311
                32'b10011110100100xxxxxxxxxxxxxxxxxx: _out=188;              //2660237312-2660499455
                32'b100111101001010xxxxxxxxxxxxxxxxx: _out=188;              //2660499456-2660630527
                32'b1001111010010110xxxxxxxxxxxxxxxx: _out=188;              //2660630528-2660696063
                32'b100111101001011100xxxxxxxxxxxxxx: _out=188;              //2660696064-2660712447
                32'b1001111010010111010xxxxxxxxxxxxx: _out=188;              //2660712448-2660720639
                32'b10011110100101110110xxxxxxxxxxxx: _out=188;              //2660720640-2660724735
                32'b100111101001011101110000xxxxxxxx: _out=188;              //2660724736-2660724991
                32'b10011110100101110111000100xxxxxx: _out=188;              //2660724992-2660725055
                32'b100111101001011101110001010000xx: _out=188;              //2660725056-2660725059
                
                32'b100111101001011101110001010001xx: _out=189;              //2660725060-2660725063
                32'b10011110100101110111000101001xxx: _out=189;              //2660725064-2660725071
                32'b1001111010010111011100010101xxxx: _out=189;              //2660725072-2660725087
                32'b100111101001011101110001011xxxxx: _out=189;              //2660725088-2660725119
                32'b1001111010010111011100011xxxxxxx: _out=189;              //2660725120-2660725247
                32'b10011110100101110111001xxxxxxxxx: _out=189;              //2660725248-2660725759
                32'b1001111010010111011101xxxxxxxxxx: _out=189;              //2660725760-2660726783
                32'b100111101001011101111xxxxxxxxxxx: _out=189;              //2660726784-2660728831
                32'b10011110100101111xxxxxxxxxxxxxxx: _out=189;              //2660728832-2660761599
                32'b1001111010011xxxxxxxxxxxxxxxxxxx: _out=189;              //2660761600-2661285887
                32'b10011110101xxxxxxxxxxxxxxxxxxxxx: _out=189;              //2661285888-2663383039
                32'b1001111011xxxxxxxxxxxxxxxxxxxxxx: _out=189;              //2663383040-2667577343
                32'b10011111xxxxxxxxxxxxxxxxxxxxxxxx: _out=189;              //2667577344-2684354559
                32'b1010xxxxxxxxxxxxxxxxxxxxxxxxxxxx: _out=189;              //2684354560-2952790015
                32'b10110000xxxxxxxxxxxxxxxxxxxxxxxx: _out=189;              //2952790016-2969567231
                32'b101100010xxxxxxxxxxxxxxxxxxxxxxx: _out=189;              //2969567232-2977955839
                32'b1011000110xxxxxxxxxxxxxxxxxxxxxx: _out=189;              //2977955840-2982150143
                32'b10110001110xxxxxxxxxxxxxxxxxxxxx: _out=189;              //2982150144-2984247295
                32'b101100011110xxxxxxxxxxxxxxxxxxxx: _out=189;              //2984247296-2985295871
                32'b1011000111110000xxxxxxxxxxxxxxxx: _out=189;              //2985295872-2985361407
                32'b101100011111000100xxxxxxxxxxxxxx: _out=189;              //2985361408-2985377791
                32'b10110001111100010100xxxxxxxxxxxx: _out=189;              //2985377792-2985381887
                32'b10110001111100010101000xxxxxxxxx: _out=189;              //2985381888-2985382399
                32'b1011000111110001010100100xxxxxxx: _out=189;              //2985382400-2985382527
                32'b10110001111100010101001010xxxxxx: _out=189;              //2985382528-2985382591
                32'b1011000111110001010100101100xxxx: _out=189;              //2985382592-2985382607
                32'b10110001111100010101001011010xxx: _out=189;              //2985382608-2985382615
                32'b1011000111110001010100101101100x: _out=189;              //2985382616-2985382617
                32'b10110001111100010101001011011010: _out=189;              //2985382618
                
                default: _out=190;
            
            endcase
        
        end
        else 
        _out=190;
    end
endmodule
