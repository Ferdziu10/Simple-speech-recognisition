module top_ssr(



    
)