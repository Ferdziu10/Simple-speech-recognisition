module top_fft_tb;

    // Testbench signals
    reg clk;
    reg rst;
    logic [11:0] imag [0:255];
    logic [11:0] real_out [0:255];
    logic done;
    logic signed [11:0] test_in [0:255] = {-95, 1769, -559, -187, -457, -200, -75, -187, 1029, 164, -385, -917, 1761, -517, 1756, 1354, 903, -1009, 1190, -986, 1173, -1951, 904, -207, 1071, -1706, 1156, -1614, -2033, 152, 1511, -1618, -1597, 656, -1084, 1690, -1733, -1547, 1307, 1058, -1872, -1737, 1227, 745, -1560, 1961, -430, 1992, 1487, -1091, 726, 1699, 1569, 514, -91, 473, 293, -1169, -829, -1892, -1684, -1279, -1674, 1655, 610, -976, -1294, 147, -1565, 434, 1557, -1486, -291, -771, 1596, -167, 484, -315, -1686, 1028, -270, -937, -130, -131, 1973, 1078, -295, -127, -684, -1129, -1964, 1209, -479, -1137, -283, -273, -1345, 1650, 536, -1928, -1484, 1136, 768, -1167, 955, 1236, 273, -247, -1256, -1906, 192, -1175, -1457, 327, 312, -568, 1753, -1612, 513, 1593, -219, 1170, 1055, 1693, 623, -479, 1862, -470, 49, 1639, 552, -34, -84, -521, 751, 549, 991, 1910, 336, 30, 945, 1421, -1119, 669, -1131, 1336, 45, 1913, 1962, 33, -2, 641, -644, -521, 1487, 1540, -1850, -1099, 151, -47, -1531, -1167, 173, 716, -2028, 1313, -1276, 787, -1671, -2002, 909, -1633, -481, 1199, -383, -557, -307, -121, -691, -697, -1570, -1518, 265, -393, -13, -1110, -960, -1130, -309, -1535, 739, 938, -1927, -727, -1641, -864, 1150, 2023, 1729, 2025, -566, -1524, 470, -1483, -145, 1620, 812, -683, -56, 71, 1359, 1866, 1979, 1743, -1563, 525, -979, 780, 483, 994, 372, 1519, -470, 2018, 1929, 1666, -1036, -428, 1173, -1222, 1021, -1646, 1725, -1327, 956, 414, -1522, 774, -511, -202, 621, -151, 1882, -1570, 1130, -1990, 290, 852, 1704, 1985, 1036, -1068, 1583, 1259, 135, 1345};
    // Instantiate the top_fft module
    top_fft uut (
        .clk(clk),
        .rst(rst),
        .frame_in(test_in),
        .fft_imag_out(imag),
        .fft_real_out(real_out),
        .fft_done(done)
    );

    // Clock generation
    always #5 clk = ~clk; // 100 MHz clock

    // Load data from file and feed to DUT
    initial begin
        
        // Initialize
        clk = 0;
        rst = 1;

        // Reset pulse
        #10 rst = 0;
        #10 rst = 1;
        rst = 0;

        #1000
    

    // Capture and display the processed data
    for (int j = 0; j < 256; j++) begin
        $display("test_in[%0d]: %0d", j, test_in[j]);
        $display("imag[%0d]: %0d", j, imag[j]);
        $display("real_out[%0d]: %0d", j, real_out[j]);
    end
    // End the simulation
    $stop;
    end

endmodule
