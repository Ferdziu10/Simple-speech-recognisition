package nn_parameters;
//parameters for dense 1
localparam IN_SIZE_1 = 26;
localparam OUT_SIZE_1 = 64;

//parameters for dense 2
localparam IN_SIZE_2 = 64;
localparam OUT_SIZE_2 = 32;

//parameters for dense 3
localparam IN_SIZE_3 = 32;
localparam OUT_SIZE_3 = 3;

endpackage