//////////////////////////////////////////////////////////////////////////////
// Testbench for top_ssr module
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps

module top_ssr_tb;

//------------------------------------------------------------------------------
// Local variables
//------------------------------------------------------------------------------

logic clk;
logic rst;
logic but;
wire scl;
wire sda;
logic led0;

//------------------------------------------------------------------------------
// Clock generation
//------------------------------------------------------------------------------

always #5 clk = ~clk;  // 100 MHz clock

//------------------------------------------------------------------------------
// DUT instantiation
//------------------------------------------------------------------------------

top_ssr uut (
    .clk(clk),
    .rst(rst),
    .but(but),
    .scl(scl),
    .sda(sda),
    .led0(led0)
);

//------------------------------------------------------------------------------
// Testbench sequence
//------------------------------------------------------------------------------

initial begin
    // Initialize signals
    clk = 0;
    rst = 1;
    but = 0;
    led0 = 0;


    #10;
    rst = 0;


    // Simulate button press
    #20;
    but = 1;
    #10;
    but = 0;

    // Wait for some time to observe behavior
    #100;

    // End simulation
    $finish;
end

endmodule
